// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Z8gaCgdP22/8xEfTb4IhM4QyAQ1EX7ngLSMVqDSbXl8VsdFWaBzGzahu+BTiiqp7
LfQJ/jfvbRJzE+MbvPB1SX1YSm9Ihd8smOnDVyyLqBxUe5m4cWSdtKqpZTfhAWBf
9BtLMFVBb6VFPyFdqAZLex0pZYZKmeu2ivZzJJuIZ3w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
Hhe5BWmgf1pC4MhKT6zT53hQCCXvMJXs7tNQgRAvRxOKvt0cQDHRXd4TCIHPGVfX
BhVTKD3eQF6Xw/VxoHdFaLPpcXGDR/vaHIkDH6WhdgS4yrLy12WMFCJnHEx4Dr33
2fNCCTBUUG3yIR1c26gPU52FiZCdurs6b2QDZp809hWpd4VTJo7LFgMDs/aiMOav
bjFJv5+9/64Z6D1MQ7E7XPHLCwSQJHwQUu9enkaQ76UR1qakHGK/UCCKKg4fo4W+
MLyJWYDL7jnlhJhEhR2xpX9edubinTBCHMOJjB9HL4Mw6Pwro1AdydnM8dKYpyqy
poxsL27XalIBRtHrmLO5BR/ehNzU4YrJk0yrbR+LW46xXz+oK/rCio4E55rLE2n1
MKj8D+b9U3KFPaW0PdFx1udfCnDMLPD9QzbaP+39ZRy5e/wnqocs7f4y70fKPQWY
Ho54xM9s4TL44q+TIFBBZpErnS8zl2BwbW9BhBSfOqKMOHvQIYcTND88IGQq6fjy
w3qGOrsVxkVOx1nZrn/Qa4kdTbyaaDOGvBzV/Rb20AAP6KAlj5Tp0Qm0u0VoliNj
ZKROMxRIMyRkVPWWDMgxMpUGl1Jmw5szIlGmaB++BPzncRoJJj2JNrCIKmsQIuL7
+Kw1Yjbww2sktLHL+mVARCzWUVtKiislD94bO7ThqE1PoygTmSzdyBCss30wLE9G
mTlsypVgypkAbtlExf5VSjZwcqsqZeDbJEVOO3QeU6w1aV9xNWnBywpogbjft6Q6
F+gvkm+HlemtstFfwbu9RPfs5d5FaDxrT/BgXIuVbTNV3BT+5u3Z769zMqiCwSJq
F7NcuPpCG1CFgs1Ln/eFa0s3JeUiJBFI+vNxCYTzZmHvKpDOUOdS87PjsAKdgjp8
HSQ6gY6w0IspGc7UVRzKPAZCWND5iyTGNC0Qt9nGfIX71BQGU23FG+opMGwHMeMI
ha2vw6r1gnte8KmHBUYC2On88ZwL4Iq+n/KT9l3/ChTEmIb1R1K8vw6lVZy5J+H+
970j/Wc5CF4PKuq5TrLSi7lsNzk2Iqhl3+1049XfRosyVpNFBmG1mVRQv98levSJ
nWSjAhzNXl0lZ/hYBnYspEd8rzx5zNVndINhMyPFNwnfxSv+2b9Sp3lbviS4qUme
6+BiBwLd4L3Kg3j/D4sW1gTLGJ8vqNlJU0YKOyB1HclCxF+GRZBJ+JVw1twfutbm
5Ptu244sg9+QQaAgyc4tCgUlonn6Crvu0+Eu6SJUWrFUiT9O8KDr9kBm9ogAXjq7
XOzya2AFQ62ml5U/fX67H6+5h8oZmxYKl6eHuX85DqUCn8MN4+UvybDQZi3EzZpY
1oP5PfYnIanaW0UfmBt++LxT4KbCzvKlgn9Irkxk6tj9OnvDh7pBjpKAhVJPo9sa
ySFcY3cZGBUMWKkZYhlGCicP2IlKw8Ic92fXSgldSoH/p78xQ15Tsmv6GEpmnest
cifo+V5yN8Ss+15A+yy7MStP7W9xXw0iL1L1oxeVoRLKan1ixiUSBRvFo7ZtS7Bo
JATrNlfKVTOwYgB/557mz1kzhItZuPjC07GKNFV+DhqQQrPKx76hUupAkZC8nxO4
kNQYh8yQJYwmw8S+R/hzup8vBN08PeSKyx0fgS6ZHXcfSysXPzAOi/GboJZTGbw1
tw9Iw7mEAbf3oZOEkk0GLigRCum58z8kEn2HnbB1ilcNyIvwpwDLUeS55Pugz9uz
DE4uhaACFA7HQ1qqSDZRro2wueKHeOksFmhCy87ZrviZ+USX1cLbKO58yfj5rE6M
GMXSnUw72jkGQsQng+mPhFRuHdkeYl8M/J3uOhBbAavMLFoBhmBJiL4PjqvOn37c
vcoj5MTyMZZUAkqMUHtxD8r6kwJY6+lo9S1xk0tpVvccZ4Kw7ah0+05Kwpwlognp
rgH9aqZGqQrylNBLKVCZQtpR+12cuPc+RaIaowWq1iSGxeNAAIv/ch4OmetQdPOK
yIQ0Pf6tzb0ONXq2Gla4MFYwl2m7m96bigChNGU+A2YtBEvYHEU7SLzU+oca7feq
oDYFiztm6aKZQ93IyhAUMl3aulkgkQZdUkl4wGNUEWetjsRhNEAG+UAgElCuW8qm
8I5lYsdx/7GPTkN742X0E+1eAZGMOLguMNZ9nbxqvGHqu0PXOFjX+XoYz8HNvE99
GHuGVAAPKplWjqJ6WjKAUVeC8otlqhUX0rEypH2Uixq9e2QiGt+qCe6vynE0DjcS
OWhHUkuCPZhHE7czz8k6qUXBdH/MICTUHaeYL+W5wESz7ldTlQ6uKHbTCX2llckq
1wc64zpkAmT3E/Wt6gPAtranv7XBt2ssVurmZ0PCRsVJwBrfjLbmXYUYHjCjzMcq
rrG54YKeQA9mS2LpMg59EjbKZv1ZQjQAl3FllSfa7tVCDZxKixEWASIaY9hKLQ/A
3ISONJL3lhx+7oAcfisQfhxI5sRs9IpdmIttvgfZubC3GuQ4Y6hMZwhZda03Gju8
bGx7/NHpEUJ4nFkVIB2fZsEpPVN2JVz1Q/zOMFOKrlYtWvuffuTHNQ43EFqK3p3Z
bLV2yceK7jfvCEyEMKa/ramm4CBoWEOIsqZ9x8jtK+21KoA02e9sa/ycoArRlPf5
ukaruF2Iou2hEgbZ8BWZf9U31GthoM2bytq671wcr1ICBgHkt4gf4+9aOqsbKJVA
dDY3ehsOPSe4My4ryRMrTAddeuVlojO75+xJ7n/J5qJwofkad2mYe22ShdwQKTp8
sdVJ0Rj2okMri+8PIAglYymMXj7ONcXKAi/6vuxCL2Hen+upbYluzwB0unUEVY26
mD4bJG/m5bvtwS9ejCvZ4xYuowL412PEQRICWZOicKgjJl3ZJIi698nynVs2y31t
SxD31r8gbfFnj1NybT+PYKSBptCg1KQ/63c5IvF+gYgBjkgTr7wwiYVg98Fg+xRe
T1VLkhE8cEjq5j9vzHmvypbTo6bMHqVBIt8GpkcM9E/aESYHWv2dVZzR75OzUd7E
aiKz4Ro10QHhIyFRstH4F1019YKZUJMzj065y8VJRfOnHx/bqrbHIpKegrVk3Pli
DgDGOMwLybFpxgV3yYd8NQueHLMBlFYyFBcTtWylfKhlfYDmm/nUaNGofln9H3d2
nQ6BYOP1JbNGxWMC/o2RvBoZawQMnR7lZMwxNVZL1f4+MpdTec9CU15gpKP2lnOn
eqOdSEE7nOTdVprfrVmREQlQYuQT3y56hTT4tDxSyy3TMiNX7vyICzKZZ/XptqHc
3CXV6vMJkpykXjUcRHFfwkJ/g3GQJp9jOa/1zzbLmEB3trskubLPJV1+HJuSVPJZ
UedoE3VaCPmjf+F3/3+BdL4j6eABbV47k94uazztCF206xKwSNtLDrMKw60wm6KX
UUufNqzvIi1i4sQDhoz0QJPN6yYFjqsVn4pw3AjHd9VVeJzoFfaoUl9cCb3ey8lt
korCHX6ikqCXXEN8Ra4NhGjsaTnukKBveaPZDSWX02Chb3TRfvIN1K9jYXC0wwQs
aDeeMlrkDyNmLl5jOu5+5HZfAHNI7CaeRMvIMqkLBcF0vWbe9vMR2mmfLj6kSWRW
8kjA0uDdq5X8UhgNDXWmhIVPXI6DfEj7buZMGwCPCtUIGNAM0cAjgHLBxv/2f0Lq
9FNTzQdEFDXK/uPzPCZ6fyX7X/T764UaMueoAMoR+27T1jsfWk7ygX+tcd2NHPH5
tj4nkQ9CAJcCJBcfA62HVcaBNQ0j+URPeN+ZC8c8D7C2ifyhPs/ZUE4jeZ0/9pli
wOTBgMAJfwnBJ/v2d3JRcmJmUsz8hOgK8Hkhlt/0FmvSlUBYRhmLwdXJ3p2uyIfC
E6qTkMR4wUbya1+4JG0sO16F8e8wOnTNq6vaie3BIgAqbDUyQHIJYkEo+b1oNdVl
a6YfiU8E5i0iaeMqTtzGfhmt5OPgb5iFMM7AC/9fXPDJIrSgY5Rr9uVOf036/Tbb
Q/z0hjdBuX21F+9JgY5Yd9Ua5C7c4JY07g58Zs2E7TFDbYpzeEKx+JzFAaJ1T41Z
xWxFfHs5hZOQsKFs2QW1EA==
`pragma protect end_protected
