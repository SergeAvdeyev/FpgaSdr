
module SFL_Flash (
	noe_in);	

	input		noe_in;
endmodule
