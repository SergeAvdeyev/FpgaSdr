-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hp6btIfOPKERYYvK8L6vJMacld7scs0P983NmXsAHCaS+n3TujKHGzncH/Dk4iUO5FzgEM9tc5AJ
lbGdJbUyEnSAayCJA4fP03iF/GmGxcmhuhuxhvYTQD4WfmuJtkXzvoyhH8Ku3QP6cEWtFYm1rel9
EzN6Evm7xJ/K+d7/OU+2xJj+lpNfnkDN3FEj59kWvfGeOilFc1sGBM7D4fknhv0/IzvxOnoJcUSh
GivYfT2Ohv3PlcEZ/y9C91DSHKA+DBxeI1SkBj2UUXTGqvmeMJ3rG2Qlo4HIV/ymV4s33AUdBUzi
bMa10AkcKHkj/LEBcN5Z+s277u0Vc+ekP+ET/g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
i0sIEIVLS7RgkgWJVXlRU5sZMF/pzWdpBpPaTnXlNOQ0Xwovh4XzLDQGmnJVRqcPU6/Qs1C7IMDX
CLsfh8+GUP4TkN7QDlQyJiUbpnee8HJryd8SAxZX5x15HUOGi4BY8ht3KXjOA0l/20dkPtTPxdoJ
3lrNAxmD8Pbpp6I7RTx4p05HLSUhgKFOvnrJctRgA9dGjnjm15Wiw26T/dLfRf/jNoGX50Ol+iKJ
qYfvqyofekvrnqMhKC6jovuWxFXNA+5LhkErKVj0oTLH5JQREnPX/JKB7KO4+uFJzmuc04YkQCbV
3S4dXtB6lJoFTQYy5Gnc1zEypQoZl2beRUfUsE7UBFgy0JVNZRXS/TSUxw7m6kQIuFfWhgrC0kSG
EhPoimGiLgmDrDKdye3SMGS49MLMFlW9fYfEnhIUyTj5+PgPtxvz3JTTDfewJpPZTpzbq78BXo+m
uBr/5j7bJTzQQyhQ2B5ndjAGef/M12hC3KW3vrhshsIO9rlMTlfM+rh8dTwNtMi8Ht6sC1Nr6nWk
Rfrz89IJZo5ah148qU1DtoWy3K0kihyaJ7HsL4cdIoeKlikX/zXifwJ+PQ1QvVubLYqaTIwFRYmb
lsB+qmNxSI2HUjaVUCngWoL3aB9Mq4lxvANMJgz3tIGZluF+os5ectCK1t+c7+qTRAPlg0YW6YDQ
WNOo5JOKXFBzgoIg6Sfi/tVHJ70XcvVkIeKrap75g2SghGl8HTakNrq9Hy79iupV74e6Pjwu1pOG
ufm4M02HB8CGSvqz9htMvwnxzyyRjDL4xHxSunSNOsaVvjKynRfke38IreTupIR2PWloi7QRcofX
fwg7lSGsPBMyB7IIlfBFBFMqup25iXqgkLqirPpanVzq/OnfNXuOvZN/XII8BILGJGyHmFgGnIMa
zVfhAxyhSlH0tzrNX5FYpOMGlHfy7ZpBRMIe8+naOOKiS8DUCe+oCPVZ7s93g8nxEtvxrAZmcUvx
m0a4JwxA2/PgICtzqkri6vmYFw3t906IXy8PPxSlbQtYS68aD7jzuln/QLF4s3KdouGQe164NuJS
xWklLE1ogB5Jt9yAi2tLqsonDwx89p+AFOHXR1yWnbroc2e1LA6lQ9xnqujCKsVMAMuJZL55Pdlo
cOFMG0EsBgntzsXbxVnQAS97IUrjcyQuU9OMl7UL12x7ajg9T3+TODF7okTqP4vzck1pWwKqQGsE
suSrsxUgybLslWdlP8Vuu30ELIaFHbmVmwErwulmixbD0HRnV1D8JZYWmYbE2MBijaW9wRKc3U2Z
qHpwpfJJgYcpUStP0abdfOojYsU/M1fvC96g8ODWRYKqqwauOSSSI2kCKoo6q3DnH9LbeU1+NjS3
EF2A0VBPaGATVZUxP2X77xNQ4UgKMqJ0esattg6thIxWUfLIHLSPqvJhxarZmbPr9vPQt+NbYnNF
CqG3Ug9OZnhoC3OwxU5V5WxL4UT57cn700R2BUnUoTAKF3UJ0bIZVhK5pfiFKNVWxMRSuBhpldEc
iIovyM70UYE+wkCoqwO+bRVFgz9hznIMoRXzw1xyqm37qkwEZr3C6hcAzmq1DraTml+3HQZT+Zeg
LYGYieUEMurKwP3WlJLlzTO+Fz9OaICuNWMrp/DM7xo7QSEU+CfGDiep1deA9zw+eiC4SaHBgSM6
YGf9qFzgVhvIthybw2YYCLJe5Tjg7Zsw1XFU3hKhSSWjN+slQQGBd+wzjxuGxudU1KHpLjgJgbHq
BjXdIkpc895HOBwZvdDXhWSHbTmLRoB0zEoa8LXID5bHbyOMlNthwx43WiaTsJXMwd8Kn8NG6NHR
HqyoihNGnq9UQbAtiLIbZ5AYWoj20FLtehwI72X6SytWywsChgzgOh1T2OAwExllAtOsjRJqerj6
+gSIg70kmYyYiN2RWsONlz1uRn4VgI+dE5nDgXoeMk6TdggcYEZUv2kKj2ojBR4AOr3FA9HGvqsg
g4dxe6zthdTHiNFAjcS1I6j8/LClfawrLiZcJ0/AfIjs7KgIFPmJQ2ZtlPFQ6587IB1DOJ0s3hYn
y6r73xTH+12Y6ds8t37LZvWyMMfiCPGL+JQxiwTPx8j+gniUz9K0NcOn3Tu7DRCbL/hQEKNsyDRd
rzHkGezxkOeZQSOXoWBlC83eMFb8JvJAdaPLDZbqDozJC53VFW0eRcjNqinBulLwAS0MWj+YFMm2
wktAW/1fGL8MK65R2g6AmxMJrvl3Bv3hACVd4wRg8gLVS0XfZ2zcsoyj9dI+PY8VVu+zvARlyp/g
ANla95G3jEKzDTDQ7FVfShNHp83PsT76k9n/WCs0D5E1RaS2hje4x9QEMXYcPfXJNMi+QEfQLbE6
kF5Vps6cizqwKx4EDxaHGaN840+gnRWEuzk3Y2vGz92VnHf71ZG26Q9rzswEqY4caQmxJzL2UZbM
LvV8moBLbX2WmG3NSItG0WUvrn4xVeruhKUWbvxvCChxeFbmdY6gadk7W9Cy/CTeouAUuoFeFHu0
JLhBXi8WyTKi3DLpE0QPK4LzpuMgLspyrDLimm1LNSa6dNwwrvEXYIXR8wSv66XRwtPkGdkJFNlv
X1OfWoLtLddpLGgyITfcWMHIfOgFfeWjhRhMySEnldsBjKqRUdzdGMSzZ1IMLjPFrfJIYaASaeGk
amJS7NNNzl+ZoMbX8EBXcZAWFugbY+TDWr8cuL//Lqm5FbJkcmro8+VhudQDQSn9vemUyV/n5O9g
xWOqwNttzkSOh29LQuFqufn1fdVCcV1sO8ZKOuhOFR187TnFACkD0pv15ofleRVMIJysSlsrJloW
TDmnRnhfDWc6FOku8ifBH2hYVYP57OyRoKqJKUdu46x0ZdB8ZkAweHBTFjWgYz45o2EKUoyfigNZ
NcIBO1XizgfiZf5D78To73IqKV2s/viNZefZa+gjiwbzJxVNJLhEs0XjQp61K/+W1NmkUPIbo8EN
jS1BfCuZZKtkWeGIqMYBzfWO+UD41z0rIsEEElX9xw6hqVmdeEhxUM0z1cm9eIpGYleOcAC31K+R
jVj7R7RuvYx3vT2WyivFbXMqhzj8ndb7okWYSzWPOgZeiQgaJmWubvuISGOnbAtAUuouDFPVUEBL
QcdWK9t66dU1pc5GGN7burcAnKZOPTWT8u3HXTD0bcMToBlEhqV/X4I3x3R1yo0eWLYM4Dxe2OXj
xGv0IfsJJKYhPta1nBrwxRZaXhJlL0V2FNHYzKr1ZuhJ54QS8mYNsKPu5inat+HfBomIahGbgAKq
G5zd+dV03A6rr9iQgSSbuqkAYSYGswy2cz4dWzqCPOxKo1S6a4kqHCQpopUKPxCihEt88Ezg7BGu
6ivpYyINI3uwY50AkL+m9x6Fb9GVYTaJy1PAlCx2zArJLPx8uQMRM63OLLh/7V+ysUnw0KBa4txv
loHQfo4S50jZD7sk6t1mWQ5fCwq/lzWK3Rs74ZQkB//3tpbqO4Z0JWbd7nJOssunl6dkTaPxc1hf
6oyigARE0RhtecTyWXxV+t3SMRFCcu3wWX4K0jR0LZb4Q8csgKhmDXyd2NBB9WyKjKW5w8qaFOmJ
YX+D549cAP+VHtOarUAQkgBh/LnWRKM9dsS0mBawMSqJ7oLnitRlxQJrhijMpFpDxM6LwSabAXVq
DSXMMFbazD+X4+eH12qVZHpwAei+6m1n5vKVyueyhb39o3Z+qVnTYKpgB4InYU70d8Mjcv/xaLcc
dTv0ewfDnlFPkU+IMAXEnGk2ka7kJfaSzpFTW2l9j9HjKTfv+dlpiUwu+mKUaDMrjohuAnFprmur
4rjlZgpOsy1PVU0aIsXi8o/BTDiOQwLrEhwVFwAwpsx5toFgy62WKUq7iuNJgfTBkGXhxxKuv9fU
rkV7m+YDqi9Izc/5fwPEyPLA7D1hTn8x/4D7KZ5Ts21V+YuyGICUsxBTK+KpMGO3Wc6wBUkSFfsZ
nZVt++j8oHc1YCxTS+hAqDToXxCCRE+6EWRGKnhHBdHzesuGQoTxUjm6g7mwzKx8fXw6CfAOJe6S
nlDaUo2YKtwK6TCpg7A7+O7enZg2pzCFiysH/guNDiXJkLKcsxXTj5gcnO3+voRNocWBIyN9GGZ3
9QFH462IH0wBkrH8xQr/tzNyVQfi/zTz3lzQn6Av1iRA8NEBOz+g6FQ3x1CjL+VcxyOkp58ub96/
fGFTvSjt6q5e+UWgxuHJbJThnCh/6/Xs3GCCiYANCB1OUeXPctMZbA/VjJ8dPuWHhSDcTM0TgTnf
6nLxQrAtpqYU9C8mAhqrSZEFirl1DZXw1wPB3uJloKkvKOEYoCdBFqwsW7IlWGJnVCUNX60kIMY5
9aICL+3NWSmOxS++ZeRUXRoeqaP5c75e5R8QHlykgFUowluBb5u+0jAi3lSgD8Uu1sW+lo56BR/7
snO7nKnP0p16YD9m3Cc7WuJMH1OCYGHlmpLNwEytSRO2jQpEXwQRKKWcXQtDdxjtumDCye5QrjoT
nwWSVOVl3TBgjziNFOf/fbBls4IVO+Z4g0Rs8qiBaV6XKzE39VvE8Yo/TWhCq313VAe6GDOaKdXZ
+mKDQG/WQsFNqrMydY53ofzixRYn6jeSCBTt6X14TcdGddolCtrv0Aj4QRuMwDsimdVqddZiX61w
OO3BS1A+XpI1IJzflRXMxSW98MnQnQwyw8k8W/bXmPfmAFnCNAR57BIp6FnYyN9v4w05LUAAIglW
EgnU2J45dp5WjbemUr/qQ0RSK88p0bIwlj0hVLWTY/+smsm8NAj13d6sLwejpq3Tq/RrSrBUYSTP
n5e3XJm8gSFL1tAwKqeg7Wd0l0MCoFZ+Kq8mcdc4LKz75YRBhI+qDMyoiaCjxB2LqF/1tYwiE+J/
bM7RDOKIXxYk6NyI/5mHlyjP7OE0+YL7OjpUk5E9phDK9RdN2fbz5e3rfDgR8ZTinmd5v1ovapSK
TcpiSA0cUuvFYUPL8RtJZgXxXjrhddwCLsCcB6Cj6beiHBfVeOEP4zYeKvez+L82yHSKiOyYlm4B
uxRgfSgVpznlTyCe0m7sCb8oimR48wuYgyPazUUn1Oi13ZhMTaxUdeecgOFrTrsRu1FW0Ztm4OUN
H4CRt83mQS0kFyhNyPTF4+funapS0JeXqkll8S8XK092X58f5L1uzcZ5Zk/WAo5jJltQcxD4JLgP
VrsqWM57EhP6CyjXNm78L47qyVag5w6//9zos8pUNcefhArN2jYigh8Pc0ZegwBV/IQ9bVXIzifu
Bfp6dl2dWI5F6T/nuN401PipMeX79mbZWGM6tbcZSwBa/Mf64zTgNajFyExeDJ0khvVNBnYc07kY
LOUPX/N/Oq3WtHHm50f7bm6biICdxHY/VGsh0KNL4cwU05Zmyp6nNwJ7VJCBcFwRrCjQ0PTzhzL0
F07ykvBT41Iov8uh24ANvCzFO7KVQNkiL7ySeWfLfDIL/lyZXAQc6EbLw0T1doT+bvajTafJ+1A9
SaXAeJwuymkEqQgdEkuVhrNF8HMRQ6ngospUDVrcbP+XC6r16XIEbT16s4FeAUZHaap4he4uujZR
Erdd2iLZll7sQ1iVv9LBA4buYJ3cm14HqH/sBEYOd1ihCycR6RCBepHFhyB84uBmknOJXD0h8oEr
eZkmdtO3ldnAH9yhwZjy2mP7rXysKdF6oEKAlUncdkKcq9w0lBT4ObgW0Xe2H8iVAOVMiWIdrEeI
9twqAzik2XjbWdvahCRjcHi2WsqZrNYRqbYqqjYNsXdnxioenpMUVuZRXBqVJdTUFIM4XXulvu1B
SnHIfMDAbMg4piuRqKtnaM1SWGLIrJnKzd/yVuKgzQt1xrDMKztXf+d80HRkN8Sl1aHR+CcuQb7d
spVenHnWutVVtKoD/xh1CCUofMokZ/DaYGM0QeLp/T0yqeVgliB5dKeOjZLOEngMsEELUgscW+uO
Gb28QtnzjClRKto+cAJUG8Jlb3WKt/J1/VBnSw0fHoi5BR/ziR1sWwO4Vcg9Q9Z/PYCjbMxQBt7L
W//mdopnGXU6Og248Bf3I6xhLLm+FLON+Klnnq2cnqCrkPugPNtga2PjLh28dDW2nE/oQ8bc3H9q
W4lfkL7qLCrIbuCl4QbrZQ3Hjvyg+4RIEqUfu//SZktXZ7tWovEntQtbaWjGu0R2rkci3ofMx9Bv
pPPanufvOHQvFgYQPwJ5gi/V4aovBG+FcmBrxHP28JawwOFuRYcVsRXBG0NeR9iPhVejDNZK5ovS
uYfOL+fKtOCbiQNm8/5iKEwK3crPCGasGrPy6aDBhxahuEnxBxSv4K/UnDdeRT+wEErE4/fjga0a
mpw9+K264KeXX8Td7g7NX4nWIgYYRO0JqPy5t4UDL/S7UhSgWa0R2ezGtvQdbDUcQt1KPffr64m0
DcsmOaGU0RvAx7RzwkllA0T2KvYt8LCg88kh/Y3GrirBeQ8W93B8SPJFonFX2SJS5jNGDxtO3SdH
HrQ52YHXwzvqE5Fo1cR7aL4aPtI7IlzeU9VQ3AH7IR7ABeeU75LaxLDcVT9paaYNe/r8N8/PgFUt
SybijeqaGnj3lN3i2r1n6Ifft07KDij5lJkp4Yk2qWP4XkUVXLy1aTskaLliFiJh6DdGrqrhIa+r
zbPRU/t9y2gbJFJpLJD4onV46OaNIdoaVlWQ9cGZYCvgAOcfHMjMz8GOtjWHW67oG7Ded8PDoxLM
2mP2BwUAifr6//Oa0JcHLPoxN3xFF0TSqNJOSuDg6x6VAmMmN78BlzME0RfE1xLDkgo2MCkcZCTx
20zTYMuXXEpJJUBBEE0bkO4utH6waV4pfBBE9FHL0l4onZozkAk4u+6g8QD5Dp0PARrbYLUyfc4w
OsfbNZXbGw9ZzE0GpqWzmFSR6WRNKb+yS5Fvwdjy8W5EUMHV16+PXoGRFOYtLWXm/9gF2yG3OmEC
l/5kvFjyv+/wF9h6H+ggsyhw5jFGBVjPnRmwEmIdFM/ffG2l71lbGzoWllF/kw0PxgNrgEm3qkI2
t7hnGRfj2UJ85YC/1oB6a1F+U+Afop7G7V7rOkcAPid5o05G9EWG+F+Yt51pRtnOhM3JEArl6oFK
8+iS3qlGcxI+tC4X76kygSsfLtxSsCR9exAjkXVE7rS8hdzOqzBVTOkaeRQ+iFRPR2FYjhxz5o3z
ou8lZAl8nryQ1Pip2Z5Jvg+RA8cEw+j4VW+t/DYLsdpMI2xScFWZZXgYAWgPzH1ZKKeftjYuSzt8
wrP356X4/MLJUXcMd8VtqV+dNFNbYjbUVxKs6uy4dtl+Lj29GJj/1Z7F154CoIgv3eFUk2PI8NZq
SyyFxOOw038u4KzfqbDmccDqNb6NxX1u5bKfavrgG2W9jNYlaA6eBzN0bIWhXORdbXkBcv/SUh4m
Zvx46Q3yD2oEo49CvT8oBZU5TRWmq4PB3jNjHRK0ETT5zcdWwEQuMlW08FuREwL5twaU+JKZOmFp
FFYLeNWyBaPnm5hC5YRzbmrirNAtWPVOqDcQyZLvg54YQey3zLQlTr5W9iJFf9m4opoI9OIj/mfu
JenlrrcHtn9FbI+zPaTDOUJDox84pnsqU8dFPLu8BCjtVzegJloW/d9zPWb1Y4EVfCPOFB7iSNex
yQXu5ax+4FfhNbL+tdV1r++g0ro9++NFO/NGQ4XHz6nodsHCrJWXQCYmUS/xm0knqM6rLnSCx736
mQcKS5vto/ajYuM5UVlfzLQU4+IAjQixt7QRo8r9QK4GjFbnm0Izujrpk7UJxXCUOdnun19W5zxi
tfE6yWsIt+y2/rY7eoZzdf9NI26/788QDlr7aVJc++t4myFQawDHgkfNFJOkV6kVX0SKWYp7nLzy
RXXQYmnt8fSZOC4KoGDalIZ2EyyWvXMOGzOL97Ui0qsaUF/Y5dRgxFAjicU2an4bLT+uvCVnboTB
GJ4d7iOcHXlpl3XqSyAgifMj8WeOUPX24kAEBS/+MP0um09KUP3A6tKOwAhev4mLF/3ORC3JqHUD
3tiyR3X/sLI/J+A/Mv5cgw89W5KAcCPSPeC2GENKvFPEu29pnKrzUFglAG0xtWR2Y4M94ZFL4U/c
7IuJf50eAEUw5MxwVyvRdAwNZGt7eFbrEywSsJ3xIyGNTkN5JSF8C+MUfpMLSWSuQtzsyELZYnrE
rD156e0XAezmzpcHHG9wbRi0v3dOvJJpNbAaq9u03K4OEZWiXzxCI7rQwf69oaBOme6cza+XJKka
W856J5G+ZGu3lHBhUw8jPn0LlyHvmxF77u3W9E4ZPxajfSRk6Oj7KwE8Iixr16DW5VSd5wUcIdXQ
cc9K26uG2dEiRbeWoFoNzpGtEsPZ1sQKEPqn5wucAOviEjXcFzuVlpW6hN1bwEB9+ac7ZTaOrvOq
vCvtyLh0jdU5nmzl5w/lROQwNRdMZ/ox7J23eMwc6SSw7Hfs3b9bUgIWKgRgO6WgmB2qUuE091QZ
uqZh+8n0ldgYPtk3HGytywaX05rH+C64sicBBGDeyEs45lPn6r0uwE6e1JwLJGTvLAgmC0Ny2Tlf
7U/x9URk8Gj2PUqdN6kI1ibV/pqvEEHi6ly0IsTwpHe7vlx4BeDfZDQD+g6cfPqXGnkyBOYvrFaP
/yP9SE6OG9dGFoxOE+Sxm5AlrsqyH19Uw/mXXAqklMVxZDMhkOAihQt462+qItQNanXJkc7tjWVr
WoxuTMD9eGeLdnRoOooxperDuQ3F6zCHXmqTQX+d3sX1ybzD0iLq/99S+KP3A30G3hWzwHlOvpXd
rUcOa/ELroIl7m2bLQeB5QYZnSW4tJ5DhZax6kA/GMAO1Gu3cgmo2PpukbWP61Gork0wb0bFitos
1cGX6bu1DAHT2K1bBA046T1w2di5UQ5jQAOB/ggSRoWdD0g2yycAl30xrXSE2RAaqTcp3FHb0iBT
+e+RpQeSo91/BjoLNOG7+Kfh37hFxQTx1uDU8AXqybby2IL+80G5tqYEn2bRRSbVzyN7MBIivz73
B4nzVPGSoH2M71GV0j9PcOxjLseVEXbeQ4vTDcXI4HewM8HyrWepRhCFYOYt6Tjbd+A8sQRDBO+P
ZqvI3rbsmxtSLy97FTtDG9a8aur/MMuKQi5RWg3tzkLHxeMeufRsN2W/0/5cYZLwB9N7IDrDwVnJ
LHPDadoMTVCDl5cxZiZ3KJaoKvT24F9qAcQkmWEJa7qjwNGNTcJZTu9A35v8wDKnUi2pcQ0N8WcA
2Dl2kJUgFJy4Pift4hBZR9EJ2PVBpNQ2mwDUCJYfYym/JQTbjdKu8b+uNzP6zcN52etUX4eO2t43
8d00tcWvNPj5wdSCaBRvXEvhKuwcZUvHVK/7CtGc0v3cdQ2HLytlB05ZkfuKQbcNb+GjtaEEXAg8
5Yhk2Mz4mbvOnOq8NmoZyEK+V9gJyjYsG0Q7eyFcRZRDwFFTPB1KGs4rxJFaPgp+TxqfHHjIpjho
UVwrobvDeF8CZNsdjNv6JYdXdQTyJt1DTMa/HyqWixRbEGMpO8KJfmPT1/kZkrHC3OleDB4bcPvl
wgb1rM4FeR50GBP+xQ7NdFYfiF0vc+vUsUQgOqvhV0id8o0Kd7pOcAKgRYl6XKP6RR/m1WAXIxW5
8/ZVQBNUsxjC5FkRXIcCnywV9hJEvQ1BHEgVPDE6sVradgx5HK7jFcXJPvSvZlf2rlw7zKZ8F15s
fpCe754pVDwjgyIsxzM7kY0R86mQd02xGYkidhtCZVT72Xul8Kk5SInuZp6vkONtld4XGXG2FwJs
3ceAe4eXThqyU5tnWw+R7Pg6PANOJLD98CKGjwx11nfqocB21vkmm9iWS0u3onpOC/O4+Ow8R1UD
JSj8IcOD6W26+wAvwF20qVsoEm+iso01iCvvi1Lx4ivLnVc3TLRg1Nzdl45e7poSh+Ywi3UyAv2D
fCzhVDHj+zC0f/uMKJ/n/J8P1vwOM3P9TFyc2FMVNBjpdiZPUX9PdeIiKyvLVuXnZu8FMup9DUuZ
bnk5O9G0lPPWlnnQsVeZ80lvcbU1blAaLWFD3WznRpDDDoHi174DeXckL9NQYfLdeRt0cC8WZu+I
sj4EAlrFG27Han8S9Rvf6f705Kq2uegiX2O/3MmtZO3+KqTG3qOYKXxiodfi9mhCN8pzTwRO/YRQ
2Krj3Hu6EyGyfGSH1HniASX/2eBAKQNALglNTkepBVf54DwFNO59Qg1UTEu0P/oUzBYTjSYpyzOB
ABV6TKFgUFWvxRH1bcKbiCxhBRVbeWhH3WvFG7Fri68z+YBV3dRBJ+Pa9rEJg8JyBObex+7Tdnme
vGb8/xLP9nxmjuTxwo0pjYoYa2i2DDw1PRpU2uTEbqdgxpqiYNtYtskN1einNBouX29z2tDVaT1a
MZLeiyLizq8Xe5NT2RiktCZ+pKDWrAmlmCEecbPr/qNwPlA7ZEBoj+x/ExqoAVQ6CNrBPFzWQlG2
GEQoXOlAjhsDhCRJxxuazOHE73fHcWOew2KRXL5P3dnfS88CQmQzDtbtZUKPnGiInNsA3Ftcr20Y
NEP8+PVUsgSK7WczaqghgQRxQ8cfg08R50Pi4wV2Xdm4JzObYD/m118W0qFAMEZHqSpT/nHDE3sE
y+SUhqCtMP/x3Pq3/bx9TpLS+/uXAgR1NFXLUVeOfQyhtSNw06Cubhrae4rdSDAGf+/I/KlKd0q3
OJXsFsoA5zEn29cDXu2WyJ1Aobh+i+GI3rT7L8iopmnBxHKcvVw5bw2PWffwNVE6ywx3Q40V5kmH
QgJDVUpkiYVT7GA=
`protect end_protected
