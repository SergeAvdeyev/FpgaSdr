-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CxWMrvA9xx5vktYIJYV8zYguijdCn9T389YRdnEdek1fPCRIk9jKo2+H+3omB1Bh6uwLLoP4xwYV
wW+Je5o30CZuZCmGfE1Y9hKSAa9oSdmfjk+lunWd8LWfghO3WuHHO2V9yP0BTDGPX6FFypwY3nCZ
rFqOkkge9rLzr3rYVz38GJpLu6ZPjweje29XamA4Gt1EbMOnUdwJkm/e/4B72RJrX54/JpNz6pP8
UZeHbCupbJSnsB+iw5CMf6+pIDo8JO6jjKhh25bG8BJ1l9OwxZA6BMEdzWJoA1uahwN5V4gND/RJ
Z53sYITDtTu9qu6G8CSW0Jv0hg200tic/LGvVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
IGQhAtkeddDtnKmjlGlCGDfgpG5emxh5DpDeLfzkGuADef5Z6E0GktepdkiPkE0a984rTU+Wj8zA
aNmp4cQheUkVEGcBOMdMcaKdRjT3ygoEDAUOnCSzDBG0VAcRIr8hWR8QO0KqH8EsbQ3niK8hwjqC
p6lAWvQ5dyZFcXGlbAYaMbIfRI/6dwHcFwcuy2+s/sRh305jo63ee+D2Z99oeK9EDUoOuDpXlRnu
uhscGdIXa1CpOmZTFhdwtTXG4Uvf0n4Y93o0kP/0HkClbX3EDm0lS0TUJl7r9QotQzpiVu99vxIN
TkP8EbvpQG5JBxMLXexT3xikFDC1iNaH9GnWZq5oN44e+ls5owdcNqaY0N/DDYRE84+FJZOQZmsL
f1uxRzpHDz6JTyGZImZSEx7Av0TqK2x7CqiFvjFu8//IQ4KBWX9f5B38NjryIb6INLn5qp+cyRGO
htfRSCcnGtDHAk4xyufqjYfujv3PFIXcvKPEWMH5NwsyS8ERTfg1T2YcMoUxiidji3QL3OeGRRgm
nYifXjIXfkAgov0RHxnwEAKHy6oYvWp9YnIgOYs9DHLht5P5jqkRFjc5/qgDvVpr3W0mjwoOF2EB
5O7e6AP1xzEnkP+gq9CVQZw9e/dKj8i7ZQkk3ka4mFYBHtVzcpnjkvyLA2NON8LGplHrdrqHFBWY
QjykKGVsn4UtirYcdHF5bQ5tYvtn+u2FnaBoXZXUT08xiuv+KV/6O8exjcWlIXPejAG5RnGuYbk0
VtN3ZfHGFDSBDVhdDOiBXi5yPvkLKyH1T3bFDsRKKPJRNqPmgxunqJBYO2pZgWkUxg5fKOhmzSKs
LBUjQkRDGSzbunNG52jQk/jtmdwoye6R7X96BlGcR8La68UvHZ2CwrVMZUCLhUHLo8yTkxsDvY8h
sFpP8TRSf78HUSG8a6ouxW6yF7Tu6eHiclFlxbSftPQw5Dw68Po9shW5jJUAtXlNk/QMJOdGhykl
QaGshC4tN1kkc8edhOdZRGnmfRYpmGR5TP8b/RMsKjOysUmUtZ9d4R7/WyruhzCPvA6MqzGhlbLk
SslZmFG1vCjpigOnYloY7MMIeNJuARKLFQh9IkP5xg51Kom697Oc0oaOJe0CPtwrrpMgZ6QUIjpY
4Z0VFh8l3POpAppjZG3BbxGjAJb9k8K+uWyC3iCUi06yiaQ1msVGT55kqVpuPfTn5sNyVr1WKsOD
Qo6QlPM1ceTBUClTy/SFSoQEUTmBxKuMHzieQRUPrQu8ppLawUjbmIY+urdhKlBNUh5ogxNgxe0F
KqUnykDKyJi27s5BTtC6Qo5brS5etUMKtSjhbqeDR/i71ekTi7VATTyylcxgNRLyj3GsaKeP4Y9d
TlgBu6quACO4A6Drn++x+qxwvACkoy0njdOoiNG0FhCG9XMKpiJkZX222tMdMMvt+hvGnVEVuAB4
Rtj7FXuCHhPj0qxqjYY7JwMtiI2EnzKbrtzA/goe6i8wWaj5oMDxzyzhcJfigC2C8EMBE5JTP4Nq
pnBHqkzZut0zvL1wgDCie8znAbmys59EJ3sB3fQlbCORG0UqgFQz7X0BLam62EzmCxXIpDWm+gjI
++lMwe9xgqg5ZQuYmzBXOGM/Q2BPVzXYIhXbtrOmXNgaf199AGXhpcVoOOQOTrdl3hIaW+V6+HmC
5TWhkrVVQO2X0gGyv+hIukK0qfTHbyLn4cAv7VNNQxW+CKomSa/mItmviNOneE5Fj7EfOAOWiKq1
TeKaGOVuhAFb7PhOwT31Is96LFCXDMWJOp+50/+hawXSl4ubFdbX/a593HALjH9/fqw1sVrxmCLb
4o7M2A7i0D4dJP6ypF8Cl03VzuANuWkhzRVrsoB7LUGnJrDTpam0fSmKvwQY4Ic6OL4KpTJZR1Wr
6xYvhubIdMClKN/k8LqdfiMTLG08hw4o8Hrt4//gDESZGPA1goEWUJipYRXyM2Dde7q/IRrtsjsL
ZjtXiJu4UbuCtNo/IJ+NUsdk3RxghiBuRSqny89hELmouhRZuxQjwiWgbHWw229Llo88XHSfgYt0
kvEkSwQSSeSolhZhWpb6AJJiwiHhJ7EcE/jY1YrRMFsDePJHED8qXeQLHh++CMpVnvqg1dWRu5RN
j/6z0c9tKXKEcKeB4PHZMoXlGVw04Ucqv7BZKbI8pObQ6qFqIpYyeNozAK944RybWY72BOvel1U3
4qW+FyE/jtZPDjywE9Ym1K9kEpId+FNaCQcsF7KtGoojDbn4qq8FUs/yip4ZaWE7ab7lj34PAgTA
hJ3McwEHidbMnLArnZULR/MKH6L77g84BbKJW82L5N4D+PizkpnBrfJgrmoDP0KSOmpfDf9372gG
tV2GYEUlAHPD/degoZ8HvBx3PdqYKH1/QNu/Jvt4y7pz1gbvLphEiQbRwmOK0Ij5A8i7bIqrTmlr
snmHDJe739Z6LNCXg3dpMUgIeQaBKuMi0UlMQ2NdVfIYqX2SMLDg0mvKHx1Nvohw9YIayhg/hYLZ
Ol00iEQN9dFlsR5lMyDPmVjJcT6qnUDtmHWRrwrhJhCCDmFJo/sL7TRmy9LCLMEiPZzqXiadRuGL
I98qiB2RVVU4Zyv5T8p30DAncV7iH2qXALLVK0Hz/KT1xYG59NWacry5sWAB37YS916iYknjwAsS
/wF9hb46p2doo+wjcePaGJ9hUFsmdDmF5qLKzvZ7OMdkNazDIJUgrIu9f9G0EwQMBXHQmuJzOi5Q
HILdY9WDMxevZ80qKGe0oVn9p2zGmO3n4NMRpuDrVj456kHKSKuI/sDNSin+czOKuj3RYFycKlbC
7stUBHuZAkgslcy2BLseKqrjQAwMMzxBpSmDQ0NimcHbXF5gY2g2TqHivKt7pNqKwgZm4s969oI7
dHmBLMRx2bniR0CttrqRIj/QqmwED4Z/1pZWy0zTf9MnSCwABixiidhvyu6ogt3IHGXrXxYH9uno
DwYxF5HkiqiDggVdoyFCG42gds2JYcnZ0CiFM7bJ4cWpJCLQDyXZxr0oP2v88u6wy/LWJF/LDfkK
QAjGL5fQhxZXJCDsQfIhlN1G72k7ixFY9V6wLFsaIN4jTSZ4ZTAfSA7T0QJ2e/r+60yDhdYsgczI
w9U7liGIosP1ZKvLjDE04HBrnNyd8vHCnCm7QpjpMdfhOv44/IRS6IYKOTASD2/bzolaqoGoRbxo
PzZycTS1ZOkLQcLgZFTmyx62OmLKShCbJ8rCsZBv7jzi2/CeEsYFj+KKeMwMxPaVnOTOuGiic9Rs
1COJXJYK0zoMeYlReoknAXzy3al6dOYpgLhhFRgVsLJ+6JBXZPbVbVZxjh5TcHCnW5u/TYkNrlHF
GNczmxX28QYnjZFEoLFl5FRtanJG8w0ObpnR5c2r+BncaNkjbwWQhgJPX0klwVSSYChNA+ToCzUF
KOGCIGftt35UNf2cT274P+1sTDMl8/JzaNPIyH9HMtw4PMIU5sqvRUaKVVeJwze9a3WmRkAhHWpM
Xgx9eiDfQMwtEiCCGhBGbYTSt+eZMNknVWricjCfKlImMjFTaHh9L537B0OL2APVjYdnqLcZtYli
+vmpFS2/Oe72MoGAGBaisHixXCiAjiqV9t61dJaWon30BvRuPo9iECBIfX0Ihyrz+/ceHQOxPlF2
y3t6CEO/NWcK4GMu8MrX3nzznuEkYmKpDyDoMdLLZOJtJnumMxY3RvQLqWBcEKCtdPGha2uUHaCC
k5KDJRQ6r0qOV3Mv9R7obIbYIOz6eNoG3450+kViMpOnq2Li6QOUbe752CXMNHgIxKjlmM2aa8qa
s4qerD/89sNRszdCIZou/oR/UKbsvfSUttM2tFl+JG2t5rznW2WQHR6dVleyeZtjVzm3uLQIT1jo
5Z5K//Dwb/DTTcZOy1+3Y2B8d27Ie9WfxpNeIdcDZrNsPkY5gn7gyFnOLegAJE3NuIww3vDnzxVD
2Fd0/bUxyKh6L3TJgCTkG2qVWyDyiA+hRJBnwHBsSb4P4g7zL+c2usg4+73JiFRGsYzZDlweCttn
DLcn4abWIJjMY203RmEuKBfcAmW8s86o1fyaONKbzwIXKZvw1nVqVylkRndqK4xxTvHRaBnC66l1
kfVx6onIKyupZX/qvAQZKXbZ+IijctdnTybJiJS6nE6nm1opZP9tICNxvLCTQQCe/mZK30dh/SOQ
fmyAtNepoSyNt8fqnOXNm2Ztx5FF0MvHpEIMHyQLcQpo8pGr2XevsQVBjI7FbiLzjpXhie1Km8vJ
VBNv/Cl2Z+vPn1wO9EFmCp3LgBYxnzIyYSojZDPPlcyoyzaKDxcJsjIW7gF2nNSx9mcPlM+XHP0t
sg/6zVNl3UdFC9QSPzZkMoWAkJa46u77v++CEtWm1OxBCpKBik67fd0otrgwd/2QfNEkA+xyUJU+
OD+JHspEtNFuElS6t+gWRn4LZoCM1oFFAIBLfvApl8iRXBlOCZLhpSNyFLRBmx5tyXvRBUwUA5J2
Wyyt037G+48Gney1IZ1PB0WnfTgLn5nOZaD17iuvugrKa9NPI9WdP3ktUZUxgwlx20Xx/nrgfPkJ
IWcrnL+zdr1WlomFRNhkfDxRHMgoI0gdfYMlMbeGWcYlEUAEqqAZmBoczEVo2WNbruKEC4KcAmrf
Un0XaAdjr2LdcdoYLYYVQiJrSWw5vFgMjJfKkZXy5kf1jHGpp1+/im1MDlu9uW+vlS7TDRKaP2E3
ehBuUdH8LparOjn1o8sJvmrPN/VpIEa6mF64WJWbbxTde6K5amhjVWprDN6h033DGvNpxoUmbPkk
ObcuruVPl1TyDq5q1JS/yooXRCiBxRs/PgdMmO9fE4Am3TMrAF5U5yoOheuxHfV38si9pFLPsskl
s7fQ+HSwoUhYIg5mYHn5VuOraxFi8VARKHdAKAcsLmPzp2tMjpofqqHwk39PTsfRCuqAuakiBrXK
AlqQVGl3muULqIIbpanPM5Lmv4lK/RiuQwDavLxGLBHrhoqHbSRVlQjg7tLaleomn6uL1gjS0yb3
dvwQ989EGxjR6oe/9p3SRldVuGtjWNcHDQ9g6TDjvtivqRcVhS91pCXVj1liI/1GYDofaQOg8NAZ
ZD2HVwt1pMf3NEjl7lNiBSp5Mt3DVDf0NTlXAxjEViL+L+AsCqkOzTKwyO9H5JT4enLV6eG/DWB0
nYp+YfVqLCTQmCQjPpoFbTuRN83mxS2OaYUQfuNm5sK3M8T3qtJ9PGcB+ZQDtGuboFcjWQ+A0mSS
pvilxenUbF3g9QBMmSwVvItKIIDodjI2lxD/Jn+rN606unfI0GNLUtfHRSM7j9OmYso/m95ztU/H
5mtViTQwocT19mHagDU3XtaZooX0lyPsZy3Kl14HKLqMHxKYewGSi5OIuRfo4tbdVTL32DHVac5W
jNK+IesEDcSCouzL6K6HUhVCkK6eAF910P40z7zo8XLyOKR4DoyMSvqLdRuATLBcO2zcOpHbzYa2
IhxNzCriq2qQq3jPhxTwcKpkZbxDjyfUM5j+cmuFrr26gdLJBreEE3XzsVsJlHWQV5yXo/tlMeRz
1PrrOqnT/A+UdL3e7Bqs5/Tnez3vZKRwdDHL+JUbO1zz6JNF/GY/Xs3JAhKHSQ0Dr08texmxxx4r
YGqJO8sH7HCMH/a89JGYxnEPO08lUPw7dClCE+pH2vVjFa4AMXXi9SPXT4XgZD0HlX0+RppWQGix
F7YM88354S0xBtr3L+va4sP9vxZBSJr1rQeD0aVStBL7b/CoB1qOfXVjygQIT1KtaEObmDnQpsC3
v6MpjiE4gAI33I/eX0HBNGkBdSzBkiFGC4OOesISJ6Oa0673u4F64sDwPnXay1LODAS03J7mYGNC
nqirjC0PJiFxQWQBmzpbTOosKIysM1SL0rDXIfuvEdmH3xiXAuhPC5fhQ8R2TdBdsHvagT0/xXWn
BO5rQdpKGJEEJnnHReHwj6krlJumlxwAg0ZGvClAHMS4slcRjMMdYOyy1oX7hpjB4YXZvy/6ahFl
yNdmJmzV6vzobis51oF4cz+N+7QPjk0XQ8fW6jzO/5Z2l5JW/O8EQ9XOW+0aIfmTbN5JLge/8s+A
/7KUd0w+B4qhGxZF9Ke6+OvgZcniWg+If/snmzyHG6t+tS6wEQs+mSEWnLhdX0I8nViT1K0FF6au
nMijc1C0OPcTJG3D/FkfooNMru08DJgZkIY7QiW51LWIIO+NH4QEOXGfQTbxdLsHQXML1Qc+8Ki5
7xmputil86YccnnMWyaJuZkhZEJxzZES09p/L4V9yxd7x9DA18wwk6voiw/+PwP0CUuM9mV633+r
/+nDP92ui1uA5KOStuSa6j2HyJZ0XbUEZ75gESEaWtBgRfMd1IP+LMpjIQg8zNVqRkE56SGZrIil
v7yevJeGAKE7FVMBR5lOhb558Uy0kCPXVmxZ/7cK+xrYp74tRSolwJFU0qTWRTD1T7tphfsHQ53o
wZQ3gY8rOiLYGL1JSND6Quh9CFuhrqctzaHzvzihDZjXxZqle7vCePttwwXL6cFaH34Vxg+q2NaA
45ZgFD+0wGCfn3c1TkDHiaFNVyCvGackF9QUDYZ5MA8i46RFp7TsZ2oYgRUc/sducIHDGkeOHGOJ
KYKTyZ3spqredGWgUhVPvdOs2M6XDXXRx5GW3CJilTncqODGyHCccmK4ZLDSSUGXq7Ze3YnktIHL
4ttzza5rUAkP+l2YPgNxNE/zsx/tpclkO1MXX5Xs4Luo7qWyW3X+FUCKMQgyXZdFEv64/+BbJmAC
joEK/O/C6A0SHznlNrnMornmuMDqahK6fDVX6VfF8/avY1JmuMA5hJMiG0pedpcLwiMc3gDS7Xnk
2yD+Eim2XH1WnGeZcBs5+aWngJogg/s85WwNXPHWfvb8mMKZ1rexIMbLuCrwTg51FlQg61EYC1go
jSjzXTGsu/DJU6GEslCrWm5+T5OVL60AS036XjHIdsYm2P4M/HWmchABqs+CLOFUESQ7WEhDAxVS
hiGo+W6cabGPVgTw93IFycmsTO1d8Kcm3KcnHBsF8oASOdRlxBas8M+PAmrkJ/C/aXbQZoN+2CQF
3B+gR1d5TIiXknceEswF0vJ+jg7o+OAZBy7PuIuAdk/6BW3FxSM8WFX6AJG2oB5fuvC8uecxJOvO
9K1u/am565FVWoH9RNsegbPZFfZGYKqDmA4rpMfFiap3jMfPB9T8rT7kfg/OSHSSuUeLCtkTogIp
fGSgmKMgprqOVZ8GV7InKH7JIaK47oXqU1bQH/BceU5NP/3Bh00LdhO+3Xpw6wGXZfWkjMDewD5n
hxuLd7g97QILZywQX/o79rCB2O+1txAd81eSW++oIWfEyielz8fs2//eaGuwcQKZeJKePVEoROAm
HTW54DEoNHit6sTT5Eh5op3Wr2f04LLeIDMu6mKoEpHwiKJf0koAkFzT062Z9Kmh9MOCA5lcGarY
4WKd5AaweqPj4mq/i5GupEzajM3Y+hfEDli0k3Sl08RqdmvxASEEVRv9sNxzf++Ng9XkNBvgZe8Y
JSasQO5tALFgxqW8OY95IGS53e4REx8R6FQBJxODHONKKGxrqIpVhXc1Y6IQMuy/ARZzK1vuVnCf
gWai3AjY261YN9qMTUYOrr7IUqPuOv1urrHNmsmUlJjhQJdCOwWMB6tO4hzb5Rb3N6xpDpN3wXx5
hoOEl3ikLWeNUmEeAINgpsAcULm37E5zle1ha0CzmBjorAvGWsGt0+lHWt3wj87yur/NRP9Alk40
q9odIdbe0ECifLNyakVwTzDRcJfTh/4hGrv9qrOhau5fSW9q0VwGFU/yuJLv1tOBkK7/q1SdNM/Z
T8m8nq0EWssDfHesoNVLSzifROIRE3blx5fb7mWO2uaFZlVyGIIQtHdkEwlmqt5BFEAOOTx6BcYZ
y111wEBn+HItB5iDD8wBv+vgX1MZHDRZtaXtxaolJCRdstBmBMsccEAk2PYw1ZTJf/TcDVZvAKjq
6bTmUJ/FCNrqOdv8n7kDUSOlIpHRXK3Zd1niEv0Zf72+Vjq2wVn4um4hxVpARQGzfTvnK3Yi6JfX
kbWZUvI212vKMVphuZ5eQz5sLO9hzIECMmlvpAOHQ/9y8Zzo1aUuwfo4Pzmt/N+7Ax56xNGvTnr+
yEKqkEqhPa2UhQroKBZjSUUQrYycGJVjtzjjbD6JOPTs9JSR5OXO337lGS9Kqlne4oO0TYqm2uuy
iSIyltmr27FLTkNjoL+HYnDv4MFzsaZNkEbq5KYnGbXUErVCYlkBg/vAYrPJjAxYKaaXyphjtlgH
X7v3rr20YLy170n0dGfbkFTyhrblpVegf2xTd4iVic3t5NIMFmYQlC5PNfSDh2ThL/PXC1pn0xFJ
YMQjb+1ANIO/T2YaRY3GpbU0eHbn1V9UMm0ME9HHIhmbgmH0/xdGPAPpxoE1pIkuriBf5gs64Tfu
gOhAjsBiNFz9bq5GtuxhfpDQU25MhF1PRe6yTSFcFmA0ex7z4ja/Smrt4UO6Yygc5NV4R/VlDjBd
wyA07Q4LHPVqeTs/quOFNtt3bkrbbrtyuI5Lnqq/6t4kjE4pI2x1+1TciuFsZlEJv1uALT2+d9b4
S377C7ANfYtHmSwk5cUBmY8GFCR2fKxwdyjp0PO49IzxNGjFtWD7+opK4mTyuRO3zlMLcej2Lmiq
PfXYXWG+/HB75q2xJ+esjNgXXTCjQ9K4DOA4rxfa3KJwenPEVn83hEw//xuNvrsdFxAhNNuELZk0
TdzDYsExvEb02fCxgKp3OAFNVhM1KijSgaibABIFXDGbUdS8vfsHUdjCTJyiazHcgg30Lw0B6Wqq
+hVczKDL/RBNMutlLG85lvROKa0Nr8mg0uAmxs7hyaUNZtxq3OmZXgJbH+JynUchN+WO7pClaH4A
6BVl
`protect end_protected
