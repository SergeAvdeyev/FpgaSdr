// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AFPSFcrH7DRV4bTUxxjtFMTLqr+gSZVdq52k5OR5Ti1/PRPj9BEFEwhocln8yJdqAqUnHQQTU9CQ
cq32gi4aYkRDEQFlO2zP6+IAP+jDiRmwS/jVA5BoSHRn5WtcBkDDl94Z+o2USXwU6gO2vO6njEg4
WJ3n/IJndBQGwwOvtXuDww/1Yw4SSSWAwQvKZ2peALXpB1ZDNmQaTC/aLmLkZHbsYXavlANKrp84
J9UYQOI+jd4tCPKET7QhMi4XlY8suid4gl1/A0pYtUM0D219lisqYSeyIm3t9bocAZCERVY4EKlR
h+OOYPYwNkQwIzgSecQxbArohDrXpaGyVVeuIw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3024)
X29xz6/CWTqD5GE5dT+H7YbVIkcNWeexGJnkDzRM7rhsQLKEFNJAPsBkznz3Y8OkIsXuHyr7lodA
36XY0Em2fvpWBVE2GEl8ys+hvpN1OTchlE3lTOPCNSihkDcxEGp9pYJIoajeZrBfJLSFZWBUJDxA
dav+/qk3fpBWLPyCU8YEDRC+ILkK24dSTeISKoizI3WPPPwkyFj42gZDfGbTp8dwEonUWn6EIGtv
6/K9G5cQvyPuWa7pA3Ep/pP82j8r7brs5W+gRHkje/2g52Hc+oZTs1zNdsweFWPWpNB30JPAsBZo
2pzpmY09OMWoPmugp0ZGqiF1MHw1odxrFvLgoy9lZlJEj+NF24txvyE2YyNE44phjsPPznXSOdqd
0LXA14qeW2aR412tiJfMEmQvy+YlgLxMNfCk4xOxXhWS1cxcjB6KytmdO0QfJl1c0mqOXzWEQXmT
8gJ8WbDXULAYDKBi6g36bXAqgAgsx2DPMuJrEbLjrKMESPoXlCA+3kIutgZQQUiDqCWmR51TnCAB
U/fV9EEqRrsbhnXO6cECTXeP4lY2AJt1xMsMGGoXX8JNFG+kn5j/OHlbGo0VqKZND6OAP80ItnKz
6IBQT0kq5tKAReAJMq1PH50fXP4UAbmXil2nY12ws/uPfJcRJnQRr5fxgPOAE+Uf7+sZsYRY16j7
qonSO9fl3T4rBoLPjXtqf1LsCmhHFhtdInejrPRFcQv6xbYHzS7OHsLxmz8k2Q+lKkrsbVdZbYS8
xscdx5f3obg6Rt3zDTOZv5tw9f2hXU1IEGkvKdCREr83UzJA9oYpQswt1nt0ofnG29WGwv6kzJXF
pP0V9HwYjE0c2ksQnwDO0AGzRw21EnptkX2MKbODj/VrohGPIK84UocZmfVuvix7lY8MD6nPwKjv
JaDfK/daJ4hhEnqtp8ijiXP/s7ic41RiNjgYSMIOnn2e/osp+0MOeEb2nkHVrFxPj/yj9l+/EGXd
T20vKe+oIDbDazdy+9JnF65Dg43YGqdIK6B0g1Sn645N96sknh9Df4r8cmn11mhqEHz+1AC00Ys8
YpZm1+fc1bIGixNQeGP6O8nYFh4RHJD7GQ1KFSQgpN6qdGsdH+MW2wJY7YjzHQ0iGJu7oAjvsvlH
IlcGqpZ5Mg4Smyp0IVjyv7ZTsTH51kDtCzpHEQRGtTv5MxQmtx8sOuAGLtx4Y6XygzlEfroetIF+
COPZK/TfU9H/tfD/IsEuz43xzaHhitQuxa+pcjIHjPVOvTAh4/sgPVXH6la8STrj/MMx1hJEMlia
zeTGLqzqLM9H0arQe8ie2PNZZ9e69J8Pj21oKkZJ+LWGn9idXVoLmoJ/9KLFkDu3YDWb8QYwGYV+
G5rtQ6hJI+/amWTbbjWmslD2dnx5HuaiJX6eC6112YMFKj2xqhH27UWP0EnJ5hc8MOVjbQZ+BuSS
4HDZQcMN58/1CGYPMG8N6laKN73WFEACworcctAWPU7E1C83eW7heYUo8ic2+CBqPNweOudIdJED
jFQZTcmCvb52BKgkWtpeZkqPmaeFu+6FsvJK+joMONu0qzOawu4ZHxwixKDZUYVh7YSQI3XLC7pi
572vwKFe1uvB616Ky4FXb8ZsxdJwbomttI7gjoDPxnuI9QpXoV1oaIphtTOIcNiTQCifS93MzxD6
nImMOge8lYAjrfGC+v2wJWcOY/vtHMI+Z2JaajxBcZ7ozJs3Qfzu3ct9y//8FwdxlCFcI0CWsgbw
CxGLv+P3pKLNe56JwtCCletXqf1bqe/iN3FJQlJmKNDtd9AfDN25VYgIec2Us/iBUIUyTyVNpImU
6K8OLXlggoy7neVuHfwkLb5YWgtCMzjzScSqrN+8jfY+5E+IIQEZucI9gf8KMNquQPtv5u0iwUuC
yAYAisx8ddWVtAfDSbJZvcA6HZ0qe1CErRMYYWVUHliTq9+BrX9slvTUbzKbLmfTJDBb1KZQU71L
u3afx4s0FOnnU0C0eSsFCnt9Qp2YzDY05bC0ubaj9JOfToZqdRQDmWHy50l17jNBU2NXfLC8H5hJ
p06NQWHrAkNU/H/5EDryPMEb2u8AFoDWjGQLOmGngHsS1Q1ZcRDYkLkz/00JPc+jM0zeDl0xI+y4
CM0szQf6dP2oQ2Nfn7/lQRAOtdLjHJZMO+W7y0Jab1VOkAzBCqeewzdViYApEnrXdktJYYs5gP0a
B3LJPn4xZrfARR1H9eIUZF5jcIfuSXO6ExWrAfzBhL5I3Zmxgq0q1fYXCC+GTrJfGvrWuhW1tgA5
k5+uufOXWbObPfrh7JH31eWk0BV8hX1PophUjli/Pj6I7B6meIUUIyL+JJdRog1FrZNRqrY0OUM0
CTWgiF3QegV3AI2Yry8wqsmzluQia9J6Z5nHtTvsSPenMbyEk8v7exMX+LgLaGaFp9P2H+SWebgN
ZHLk1C+mH6bFCUEP35O2qK36uM6w/OcIjkBB1UXw4Dz07ob4ZYfv4lBPsHUqrg9qiGg5Xoi48kWw
FCt0HFB80wuMuwFhwfw4PX6OOK/CgTA8haqFB+xNUm9JIQjq9N4kNlXQ2aVMfnhlU7+T7Q4YMc+S
AgHnA2TVIrsLc/BJcxo8gx1RbDLQvpGQgZG9PSX4njp85XG7MuwKXyPJvpdCWbCnEl1i6rP0bE8A
sV1iD64nSliMuaRM9ENlx6ue16PIGMAUpwTZFOB+0Tponlb7BxCl06R7Pb/PWpxtbIr6+JOZZLwn
+ulAer0YOl/Nrv45bZHrtJ1B7UeRONlpnPa8cDE1IdrZ8KUGvT4I36L/hb0aOo852sbjf3dO79Az
JpyTLqerCmIo2JIRgR6SEUdzFO68QLsDg8IBh3IBQpLYlxKA6veX2A6DgnsGzidmhUuwnMfiyvu1
N1zanWpJ4C96lsfjGYZBMfgN2XFRw4hHIvhAnDIPKVNRkgtYHwzmExl/ZwC4kPScti2biYlUFel1
E/DDgGF7g36ZRl+O8F327N+jCrvt0gSfkUSS9EzrolURuYB0+/K6UiXghQ5yTcgnioTSfxVOzNOX
/PImkX7MUVkxIjw8Pj2h1sTQK0yDLhp3Jv87iXToo8cNbyU8szxNEeaqvpn/uyObvluYNMJFT3cx
4xlInb2+zS5aTyQDdyhE9T4YbSD2OmyxvjSRF3wLwQ0ykMbMfFNiApHDvAoWvCyzCX3snRr4eWPB
Gkcays7uOClS+7Snkh+FSApKOvzwQUbLO/oc2DEt91EaHLpsxlNmSisrRROOCKMps3nesMk0J3bs
pWWFUitv+X4TqIYTqeNq2fBaksLecccrZNrioLFUBDZc1GQXgVX5J82CrK8yN4QzycP91dmo8eM6
29qNQv7dkc18e6M3NxsklBJb1yayG6EEaXR0zi42cJQtfU5jStmcfl5z9J5dSGPF7OTv++AZG8qP
KUHqYVGU6/3IMr0iBziJ/fK31TZq6O9YKFHVQAhUw5sD7UKgX0o+YWgktNUJIIlosLMVU5maDRY/
EdbVDUkX2d1q6KqGpIFf9hw6AfNpk7tKqHVUDdzvSLJB/lHicls4LylJzFSrkESnvWQa4CizFXWD
E16Y07xBVEid+1zRQjOaHS63O4LtKcN3ebP4ukikAqq3ShlC+bpKxBsC/u1i5FTD1ON1OgGZgUI1
q/emSW2zz6iQw3co4mPNgbeePocuijCj8ascOkgqIv1znA5olmqvs9FKr2MjnOg7cjuUt0HHrspL
Ii6y1jOnogmUoJ4J1n23hAVKeYVlSONCFYc8Ac3k70FwEY8S0aVC/A6mnm5k0eCgTFmP+1/lq8QM
W5fh+nTL7eRY7Z6KH86/xYfJeOC3NzXxOxkbljwEjLBv3l6egecB5jcYvVNqqH+h2q5gUYRr3MTN
QaLIlYbZLXUIh85HeD3uSXUCXXLTmBGQnfFYqopHYWSTptfq2u/uNaR/I5in4tSVCvB7uiiVvoA1
SqYZY1pfhp8e0JFmdEWcWLbA/YVsioF3nsGVjHUxdNugGUBbLFjeKFfr3XsgeQZBDqmg7lbauyCv
vxBw
`pragma protect end_protected
