-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OyDy23y0l12To2b05k+7pTAE1X8+lcevhmZCIEpPYl9atS3qyWxmZ2kvtOSuOTOEqh5iriJvlBKr
D5yZQ/8DSUijc+F98T8HnLBx57xDkkl6apRmLoqLb6tzaKrfpsdZ2YIjwUtmHW1aZQICv/I/4eE4
zZR/kA4IDi2zUiGXjazIHH1LR0OUmw8O+CQk8NzqN/TrdIr92zxk4eLiVK4lJd4mxjfrQxo4vt+j
3T/iO1+9tZFrFcm5Kfamg5oLYGO88NnPpQEt/dW4Ng6PzgridLioYVhEl0cfyptBdwpRHDJ+Qw7W
0g/FPEhTilkz7tkgWt5df9wExpGF3gTbEe5P/Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2640)
`protect data_block
obm6pG8qmpqrOu3x57vC7aIRxfbiRpwU4NlJTpHCU4u6zT2hbC6aU3uw60DTso/hkZCR/pKGJYKP
b5mpCLzY9FR50wDr40J2/jWO/9TzV+DjuylCwM/sRZwDG04oNlQN90sJ3Mth6HxkQjATBcE85Gxp
yGh/N5eRkhU/NVI6bDS1u4DxuB5ZWZPBn1DXE9VsuQn4clsAaI6EK3BJoL0FUG3O6uM9NkvptSpy
SK3/olbHHQFry9EYx81DhrMisCb5HCIT+5pxagYf/a4oEXio+ylhY9ZAsA3d5rwl4gxkCwUqg/Sm
GCqQggI4sJoFHFJVKYTxp7gL/lxTAz137LEg2GkY2TW1U/zyJJzRRfpq9AWBPutHlqKlvIvV3SOu
MRE0Ee2j7O9hHzatYXuehJK/MaDPCJ5JUbSDg8j10G3lZVJwJ4ihzvOmA7FiAPDoYUArxviJn5Ee
a8HneQbWUc/tyDLjzOwzBWqGl2gozJ3vC9Wb8O5M+/bEAJlEwgXHv3wQkAvI+jn8U7VfuBMJA1rY
ZpZBQ3MJAtx2DwNzWYP8hCMi5buhKjPKiAfZ97ukR1B8S82/l70cgrIGDwSvlWwdtwty+rAmapPo
VzEqqQOs9VSsNy00A5lWmr+h6bSJi9OxgMd8f+3/hB68AWgzcdj3VLMx3sfU6fbk6w2ncc51axjr
b25rJ235ZgWArVr8paM95DH/dsR01zFL7XmqSYLougrTILlMcxoYnW2OBaWrjMDu1+oeq8YSAVsv
BtiMWCALxnK0Y29rdJ9SIfM/hEi6eO+0QboK+494T7bS1wmbTWryT9sWzHORgQ6oJLq0pGEOapsR
x8SnGTpt9fRYzT3lVS1r2nhy731Fgq86VKOXyBCp4GTToenLLJ1gR10A01SGjaPkc+dOlKhzbn16
1LRun4HKuYnwn+6a2U05sVnXnrNg1RHudNj0F4lv4p6UIZJphTQQYsMPr5Ef2z/p87SX6r0Jc3FM
Xe6fe7FExnhmtq/yuqo5ajRCnfLvCoZj4aDsqjRO8bqxyy8GV8nsxZqz1ach0XNUL/YjoxDJDiqh
rWaVEISn9REQWJUBuzf5QGoeqJ/0HZjn5hkCnznHOpboX2uB8J4aYevO6vzNB3+CBHdHZCz1cXIX
FypDQblet5TutKrmKLvRQNb5c3islvb2t+A0mLuQW9gznsSc+DGhOGpTHyqnjagTyPrjlPrhnU7u
rdwy5sBNOOObUweG0nDKZEOCCMnTsiTZp0XTzcyt6kozt2gLisaVHvWcOTeDM8s2+61KP0iW8Vff
Rfjk5WEIDeJc6cITa+G6RuXqEw9jdZzNpKoxMW0TwTjq34zT72eadS91KlLRf1K6XrH4yYeAqt6N
hoD5PtfBeIT/s35YhlzV40WxNvGHOs3QmX07MlVSJEVOfB3x3JaA8mRbfYSNZHgw2sWEA8toz30S
Oxv4leDnlKUpbcWgJBlpno+nXpcOkdeviofBiRMgGdOzzJnLBLFbkxTcKqhs+LQdZnvfhspvVjRF
ZF2/O5hEv5qAHaZiHZWPCE5nVe/zfG1ybon6lFmNtrYZl7pfWivmUKL9zYCChAsORi5UVFHZ7kEU
lo82pZ7KmJNQmKmE0aUeGnW1jCP7P3h52vUgeOYp557dSOFj2YzoaxTHC8U9bKXUgvTs/lNWf7VL
yQewT36mwg8zaSdfgZJyDoMPWH8+oSimQOaxiLpBu4SOqPVNFC9tj5VnHE0sBOiQnhtqT07mgGcL
O2nfYhai8YxecyHxuSmSEjTNml4D9lPH09OiqMJ3CN45mz7wm5CsknSyldkN51mCzwKXVeyZypM/
1PgC/7OYjiQnCJcqcmTnvW2VB+2BwqZX+2SIoy0+coBQN5bVWW6YjyYW4ZmVe3hvL5L/9wnlkzCf
NgfzEJGzqOiQnFzs1mQ8zwlbqW1YqlTfYBLrr+a/hkJ4mJAIGwuOrnUgX+tK4ObG5cHpCXdHY4th
E7omSsHZIIgkdk2Gg8KkmUNFRJgMs76vx7M+xdvLlX+Z3Kw/wlDIvTGnV+ITiDjqM6Z1/g4P+Gm8
sBPed/Ot4kcFe3TXosvhvSckU41y4ZsoNhyqGW3U2UeCgPzGSRx0CiNER28awkWPktuz6DM6YCnm
af6L9DmR4DVP/VscAWfKXM9cik4/X24rLukwWVIrf8fNn/0vOhNEw2NVPCTxvbuTc0ddMHUzzd9K
gf00pQzMqgki5jYhfVkM+Htk/if/rhxN5YVoj54wk538mvUqYZnFko1l7R6JtKUEZ78I6mQ/aHXA
fXbUhpjsTeDlDSKD9FstzIRxIW/ZPbhrtmFDjucNwEuxXyghsVcu6kElTXC+JKnFombryL0rkuzp
evl3DzJlqw+aIcj6NeMNosEpmaKBgVRsimnl9NC1x44RI/ox93sFkFY31AmyeKFnHbHs0X7oiYPf
+xyG/xIwfb8QwR/4NIvHTokkkk0bx6UbTOPMbFwISCVPUnwajscMPY3TjQPOCWkW/GCy3P6xX51k
i/oHAvAHy0mvLCIn4LU0X0fk8zivmqrM3YiiD4NglI1Up+YoYysKxaetojt4OLegiZzn4RXzS1gW
a9ZIAvOIdpGljT5P2mpTpE6VdMfR1aaUQK9yX5BMbkeit6ESezJ8GylNF0cKMC9bJj0Vy7MTOIQO
fnCKntBDAnZXsy0+kckaGJsi8JNBPWPIb0VeBHgeIy2OL3TFnHvTuqcp19nAsK7S7ZWuqAJW3E25
Y3mKVAPxwV22p9bhUS1HHXMYNpdFFZ7Ly7UUOnW1kdwwKR3pmvcDF7tJCcTWEqzrqQhkOtzIzC1y
YNGe5Ny5fQZnS+qfhCZnfm8s5wFeRWy2zlMKUYWis2CTRqK50FKGj9qzimUKejb4pWWxZe04sgam
Q5Mx7f3GJpKX5pAJJBz5bdivtc9jzyMaltqfzV6LyHkjnvvf5nKdm8IFtOUCca0k5s8bDY+YPleX
rIDJ4dQZYzWsAfremIJfn92rtyWJWa8ik18y4IVloFKrtRCWB+9sb6c0OlcHM9LHcM2u/u2Ky0z+
CXDQs0rdToL/scE73DdmmujJtmN82HOBTvHErITwUf2ost1JV2JI8ghOV3MhCiXGP7ZNSWHpIYYf
oy3uNyvI0lq/15lZcDpNCIMM26xggliagEEdSTeGJJmzmLpmWA0DcmIiZD3QO1CPs7JL0+nsuiId
UmdYoAxbCp+KIFQYft34p60U2U7fMC/hX5aMYdxgrVz0bwDBv02tHTsJbn0m/BQXWWOdS2JMyXy9
f2E6i6/CHIQKlr6iQLrGCabdrPEOZ4eYNXiVUskqIm0wP6jJRuwmxR3/2NtNDvi+FhBM9vYPkBnH
niLbqsAYPSPZklWtrND02wxXJ1+yrea6Ew88Lj39gkn5lV4RbwUWFYcHqgNwIn+4m3Nu+xQDWMMU
mRwBSWMPVnh02io4LUVHvxKqz8U/eR8YOhcSw2MzCel4jC4YUtNzOtJx00fUhlX/mVcPb99TcoRI
j+JKMGN9uN072IBVEwnzBj7I
`protect end_protected
