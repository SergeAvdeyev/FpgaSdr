-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HpQ02cIN9l879jQRWIwL8Ek3cGtIaF2uP35PPKxPxAD0qECV1b0ezWH6nX2j1rm6uUZk1mP4txV/
F67zRXYdhkVbEV8eJlOj5zvsd5uFzkLfkLllvHxCoEWN44SKvcftBoHYWnSlNHCSiUIRcbD5zy/y
P+hei2upH6J0Ypp8uxKEMsQCqgaAhtkazz5nS2zDN/ztECKTVGFQD9uwrgQdao/YBXGKiBmLIcE/
GoftPY/x1jgGz9Mjk3vZUAJgYQ4+OkQRPmXFf2Z7b/wKNVRk8KqdrQX/hFQTAdWuowj0H3qCAOQr
/WkCDrOnpN5s513SxPpqguTdNC3fvHIoKh1ibQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
l71iQFh2LhR/5FfvcDOj792C90ZtlzZBpy8zczuCfcVht15JcdN8kXUDtEWBhC4+/phvbh5n7JRz
gWP13eeJ3JTz7Whkzz24VuZENifHbGxsnWh5kp0mTsdbC4YTG6AWiPNLLciHQe3HWsfXkIHaaWgx
AAsE4F0VD5C1M41vZce6ofFDk3Y4dIaCmgHeTEnGN54aQckU4CPZKoaSRL84XiQkF7rtL4aVxYgW
oWFmyQSHAPy62fs+7ef0WfEHHtTQ2Sk5o+JCN2ijCp+jYnlUovF/MWqMZh3vyTw6DMmHrgVM17Hv
N99WfLVe4ho1fdHVs3UPu7WVjlpi97AU1OUNAknsbrhur0Q7dLQFbp4ca9Q90GW/+JYEJT/1A7W2
FoItmt8PoqgFuT+9WAVFYlb44/10S2HCWSqDlNV/qW7ikSn28giKAU4uUZEkJcYKVkGUcSbnQkev
NsmQgOncqGe6XDak0kE56ukqPwpd6YWIoy2PndvGFlwQDTYYNN6QOzIV10DJt9Zt4UVhLRucXlad
Y/YfI86xNZWDliT5ZndMtznFjxGUdfHDeiqn1K+Kd5cXz4QxfRVQBd9APPNt1rEAiaeorSMkseAA
jY8ItDEyO+1VVKRru2TD3Xv0hfu/gWgyfuoLLaJxL5+cZz0EhedjrKAQNXunPuumsElvlibGqqJH
3vbnDiX6fToekN3Mp5tMqxQX/WwHXxQ7kt35frDi2AgXjdH62q+kznF/yKqHGDX9924rcK220rK7
FicXcj+Iz0yfmeYar7Nqlt2gOT/GFx+K8AfthjYR5nZ/A8x/CTqldjn8Ijneths2zX0pqAjXrRSH
dUWDGOH3MzdJ0SdhvtZLgYIyAifqXGd0RlsNIL9VqVZ1sf8dpSoK73BsfyNZiHdrpCFmZGBii9NU
z59piiDbA3Sd2ZGc5XTNsEXLidaGlsXGJ9oBp1yJGWh0CDimM4+kvSJhamqz91xFByPdmRJG0IlW
MBPBSJZBXN/0UcXV2L3ohKycUmNf+UN9OE9lmwN1C4a7ALZIQYJopcQA1c/amKfsw8y48RrHG+Xq
CSnANOiSCKl0rsZj8ba8VEUYyHsLvkWTn2cI/tBfXViVV0V7jLil6sXZ1MDroodUVZmtqhfv0T9W
rM3aXX/ehHvlNwU87NcXinyo/wwHSgW0XASQnHcqJdazKwxsoNwgwLZ30vTSXeyGZR+0gZZfftRB
SR3uvNMK3necaGR/a4wuuASvDQ6Lp/dpVee9gTwZlb6lacRqRmYokiRqBzuHTJZfKSrFvJ07GFhX
cW23M7Ln6e0n7ODeikN1tzEIDGZib901iVUq3naPS8n9CJ+Q2dd07RK3Yg03w+Bdy76PFY3QL8sY
iluZ4KMidW3JOB2NTju819syONfNGGVhjmOT70OHyy/3csCIv6hsYJ+5AT5gwLy/XUKWj5gpu0dY
x86DEM/M2OH0v2MlqqJ5I7exjhSh8eEU6Ziti9Qec4HUARmnETceRMcfMwjxWG8HHk3sJd4BIeAF
42ek9vs94hBxqKWrgQQW8Gw6KbjKS3WjRaccFXPpWQUqwpG0Z1QOOdf682/5TQO8PdkvYyN07OS9
uyBW6A5BzcbGqGSqo2y8GWMe7OSiIS1wjlWNwIzlGM0ihr0iPvhWfgsXjt85ItYXO63kC93KPC8S
JKKE0JBDLeHcfrPLkU4aErbKToC+fjoE4qN8y3VW0NGE80OdGPgoFAmBmzqHvvTCWBfxe8dLiAO8
UalsP43cBG5wUlTFa969tEmFmM9Ty0tqa7T1bBPL7uMkBmX1il+3T3DebQvB2RkHKcpDSLVUPLYv
r4/YCe6JtbbMNnBprNqlTMlcy53jCdZrGWnNuZF6J8irWQfBrrBdE92XGX/2RenRoW9yB6rjMVZ2
GDgiYb5PIr1cMWbnw6UODqBP7W10g6QTK0Q1r+wo7xltd1pIFzXssJ5cNSDnCTZasDtMR0XIPmIc
RTTcNlbIBnR6Aqs144JQ86RVF8ymMeRLpI7AjcsCjpSiwnqbnVWkFqlLzsXgGh+hx1ueMIGtFl42
k1iSP12iiGWY2Er5f4xk+Zr6rLexL4RW3C+vnDaOshFFjo5z5VBGYPCfd3VGrAmfSM1lzYIuvUle
GEsSR0o1LBPcuKDrdbvqnLQmrkgYi7bO9/kybjHv59St1m80aMBLWLRiqVe+ZiACmeSqqczxZ6YR
XHtPZxuvms0WKcILdctWL0zBpcQ0wPBdgiDW9/K/92MZ3e90dD90VN0Xt7XqE/GyRplRknaKrhQ0
ObpaiyeQeqdjsKfUUUxwzDPChsytuKZtJbaUaEOdd+8OoH7d7qmTSDml5He/iGOTxQ1ZGZWEpRjY
HaGh6KyMOI8YrBV1L8f9Pwfx81rdNUk3MKak/GmVcP+36qpcIRebkSQ8C2jsHihOjF/wdaWV5DD7
gZjmthRPiA+tluOcEctKbcRZlryeBUPqrkTeE9J6c55RcxV/nrJozDazirE+N3Z6CJiwOzs7zxcw
+C0N+e30l306FJ6f4squOvN1Xny9b8mWXuE9nuAVaP5CxXcMjaTec5xd0cE3ysVeRzTIdNYPo4a0
4m+yxqkhxS1WasOsJs1PeKqW4MR5CGK8f0U05NF58I+yq2+SFcFvp9QhwZQZsd+mkZ8lm6mVxMbV
glLlD2BRA837HH8dl0J1KmMI1HSrXFj+pbx061KG8Q1T/ujcfKf1FU/PJRGNbhgsb36af59ElRSP
yyeYT/I/XAD6GbnO9yAkJsO5jfH8m6O0AO62yLg77Lm6ZoSPaNDpy7pn5YeWV37EXcOQN+0qVomZ
UUdBWy0F8fWXqFOkBAGtFs9PFBxUO17L1WY8TF6ii+Ph0j+YQRd7+gscRFvsok+R2BvTnFnOFbAP
tueA6YHNTDp5YjpJM8tGD0T/NsDAMUMcGla8769BMs/kwLpB/AD1Cvat69rVxPUBCEnciyLMXK9u
K1AK+kBOSUh08SP4F89qfLyWx8VfCys66q2QkqNWCFslcXeGYV9FRf3n8S4OaQFLXrYPnINVEp69
Fmo8zLndTHJYMnpmbwHt9CgvWIqNEq/jvmbImZqrHdqsNAGSDcJ2VhkJ6qhGrZ+0wJ8ZsDohL0iw
G30juC2IwrWb+7ZcvUcj7wwMsPlmiz6OMRghXzEdx/CS1iciKvonpOgKRr1TfIs7RGukbrwkD8il
92WtJ76cwFgTxlE2TI6xK07izIxiSTTra/zP9BJVBfDSHq4u5/ce2xc9BlVMh9s7Rf0xJg6HS1e4
tqpfLgZa3BmtkwsyYFFHWZHjTIt/AM2S/f7fMSIDb9kFVsEK1F6PTRsMGMy9m+ovildy7ercb8In
IQigWuM/gXBfvjteemjUHxB01nTVE7rKHTOhvuTmXncU5QXdCS+9uUj6ZI32WPCXUW9dDgXKXn8p
mA9JGjsASwf/1TSCa+fpTOhdPXSsZycajWO1JaqisKKPQuJQewX+JLhSp9Ofc7hKwUr+bG4n4jXB
/0RQRV/BdAw4hR7elvNMWK0YWAZrdLSBb9IyIssHFkcIgNQeWjE0KNzf9JJmo6zgbE6IS8MYft79
tGOL090SBxwVbHbWbrdA7iGwi467bLWYPlOMotAM8Av0D/YFeFtPe7LylNgy4t6n21IgmC9yBHHe
IQlqiLDzcsnx1VCS7Ipv+2HMJVOvM2yNsNyYLAc1aiHvesJOMcgXT09VZ4vs6Ggi6gCe3/r8Gl6e
JA20QgnvXQtdJX+sdflWr/9d4ROceipwDyjEp8xsfxFDtR2NW8+xJsohP8ZFQc4T6WdLQ+qD4KJg
wjbD0YCTQYJYqG6tVvC9CZkbYsifJiRx5GPP+yCYsw63DMREIHU9BqtnTJSP1wk+1xyhHIlL5eIN
KL6tNtx0kaQRw/nSXFvDuxPX8yQFTPdJIrDtN8KIN9attUj+jpo5MulHUFCFI78vY0LopJDetrk/
Fk6h8uE+EzmRGYUjD7yuW3NQ5N+mxp37NsrfMmonT13VgglfzVfOIDTg9T3FEDLI87LyoayZmy7L
c003d8nTdxePiy6B3UM6EzSSn0u+MqNcHS+vD+YwsZWQ1J70W/BoV+X1Ng/i8B/qVrsw17T2keYY
XFW/aY7wzx+OdOzFoi91Tl16gYaHcygej4JH2uyN8yIDb2nuEc/1AinjLby3JxyLrPiBYYqiQy6n
yi47heXAjoecUQo4mktICxglQUAYo13y1HpJk3KWIoLi9a19XCCBDNXagmpoUAK+UEh947rCYC5v
6MQq/7oyBA4oTLupfxhKWJAiR3BWVrGNVR7pThjbJwhugD3RPFalrL+SjSip73snLmZaqdBSX/Lx
tuD/uXLdDRZLsy9LeD+hhuJ3Y7fZiNI+VIGKrOyuFfhWUL5YvcAIkoH/C0tuTFt4tk7jiNgKlMuF
DtnGrRO8TgHu1AP/3oZ+xR/wofCaGXknNvZVLe8z6n3fCAsPEFywYbYP4Fyj55nWvrRYScrgBEyx
zbuGpUqrQ1WvEO0sTUVHwEBlZEeVsEp6rQSFKyIxwUbrgBKKm4Tf/+D18afjxrVmI/w0hhe5ACFG
WVUCbJ/UoIHyTPzDkkOu/GZvZNpjb0AvPBp7wEzw+UbZGvmU3xJzTN+W6A1OFHGh0pO8IeLjFXse
1/9L+pNLgxseBxRwc4xS2wfX59bwXeT9bfPierMjpEkJtZVlxBWuqAwYZoR2HNO8puywp4orKsYj
EJBhu8tKCCk1MDyQzz/CWd9Cz+KRQI5VIoEZAu8i6d0X5bYz9hyC+1wlc8DkfalKgBbrgQ9twHXp
ZIadRVszie1rglVg8iCUptpk/IfVcuhshff/FFfBK6ozs6ybK5vMlqE+IkC7MIizCj8QE+Aak+S4
96dzhOjwX4XTGdsb39CeMZ0lYtv2uRL+6F4mqi0vLboEcgIHL2zi+70lTaMWQkbpBExmdbs+VMY6
BaUicAOJmFsynw05B97PplDzpXkU8p0dyEjoHfVNxs2vLP6vEhIA+N4z4hR9LcwjdFurBn76iMmK
NR1On9EoxDnaviFmFkAMlIBBqt6aeiVwCDGrNzsj1rhGQCoWv55JtBmhHvc9wowaRr4RfwaJNEtg
go99SY1gLUCkr7gxYwAKO2MuTaRCcasVMr7tbBJ/F2oTZaY+uEEteO20NIGGxYB9mRfMOK1svrjw
jEACHyjtSszQByChQNC8RP3bVyp0VDn2LN3uQXMOu6v4JNm1tYqhtZ2RVjCyVO7ibjaenZHGxmPZ
79r8EshmivWFfaUKuREL1fCwab1K1E8bUjzrvop5Z0PrOmnTjyqQ5WIfbmT3DDNyMnYHVGskt9lm
eo5Poe5boTrMDHmIqkaempR+zAV3PcneOLT4cuvtMvj72REWMbRC37YtXSioRLBuxC1g/TAWj4ic
xzZk5HG6KbK6q1BWFvZnk/ICoV5i6/7rc+4buADWvbUemmYWzdZv3T18tuDsEGyZWSywHvu7MsbI
Y+tFinFaILvsm+SVf7JGMlaIrUgSG3SgT7BPn6Y0uPz5KUHIDSq5Zw5qYasYA+26BD52IHrkibPu
eZRnIxhH+gEBj6yqI0v74OMIS59fPSYQrhe6n0XVpUpva8sMhkhNXpbkF+xoiyAvtbHj/h4huPqy
jjlWVl+dPa/2PHljdHW1/L9R09gkxhz+jY72u8YYRppUznb/0ro4+ARYUgjH/Oj2AW3pwhU+ptBd
aFH2xygVGTh80aJLGNHpenfMH11rTkc5eVSLHhgXIcOt60Yn0tO2eAwnqNnTclDBbVtp5bR8V/he
cWLGEv78b8PN7gW5Ulxpe4ycOe7IEcKnhhZqKrTFK93eeUCT+0jXyQ0Dh3hJha72B43XahGalL9e
8NbZFIpvsf8wywmMdc5qO7THrItbvAfWZEcg4gdDYUjMIKzC0YRJxl1N+9BrbyJC2tcgCMrbo1s7
vf5rUd/FiiYbKzffG7P+u0yQONLmU0X9hwwxV8Mbs68NAk32XqnC7vF5gvKWjCGWMGoVuPTleQpu
BmWjdV7dJgiuIcOmTScajND8OYFrAYCiG0vUUdBruJpcy1PacCPXh8XYDzPG0d45/nfe9sHE4wcL
SJutoWw08eqsTaoXMs2agdQce1eq4kMm6geUydNLWzd+y1XyAw6eeCHp0iGjceQsohVrRdSFd4YL
J9XFEBmZ8OKSOXPTBv41D8ww0sAscfGCx6aBW+6rGIoW/tnicuzNjUFJI3v+PiA9Z2tUDU4jhrFh
QDtAW6vhS+9ydUY/3xvCOwThcCbS2SntbMeAabvZZ2WTIS/FkpzKleLDrhkiZXNrJOdZ4A6YyvYh
TMXsNHMEhZ2Hjl57yQIf2rZNTptEdavCkhPTnQxJ249BvAEwbPkLfkyZPl9peUq8zupazykQLr/i
1sesWkI+4tPEokOkHPBdpOat6paJbw1+TMsmcZUpEf4Wz7DrILCTtEAmB5MYDehpJP0bCnUPz3Ti
29SpNZBVFjHtOxUY/4UrMnn1wJCyaBOfQ4j+d2eTEI9hLL5opU/QmcdOJE46FNTDqVEpPZdgiJPy
skTmOI7+2BVYDU5xUsOxZkryv7iWjp0eiuOscCNpEmvu1KASC4Xxywk3lYSL1QQdjWj16TbGmizr
At/0h2uNNKeFHTPnGqRAP8YuBWR7ELKCThpP4QhaVBSc4Vz7uFbJNRCd0gvNhRHAL6AHp6TBtaZB
93dWTaB7PDgL12DOKbKHhRcBterOd3ZNIJYxpk5KmPg7IIMt0rfnzSI5aRCaKy0zcPQKFb3QvpUV
zLvZW4AO63SxoRdiB2Kt8Alv4VnyjAnU056loQPtO1auAa6OixInAvwI6UwPwNYBhMcwQhzcjynH
0epFyM2DIjCVESOqvzhQgn/0Scx/+pCUBpoFr3ZW+E2DAIYdGObiV7OBNUeG4EoKej7Sks6k1M5f
PiU9z5323AjJCb0Id9TGa8bX2eHrcZVc2vnt1Tm7lmuWQNhgSGGeGikEpmn+rHVpCiZjRrhYS4cI
kupgJNQyr2w+WD/4/IYAKdrQERqHvXTjsYpAAde08N/8T9Cbj6V1h0Mv2WxONqAOyEe+/LMfpP/X
DU3LngkrSMCw5Vp1HJpyR2dKS9JsnP5UpszyFY5PZco9m8rIgF6ZohswwDYuA3bqrcv1tEVnvh22
2wev9WlCl4rCaGKSl4Pj/tI+uT6A6wRj8AbozdT3tkz2AqapHxsal8WK6iMGphPMfbx89iZHS678
hmWwmYUHGQXtDyreqQLVCrqUw1CHl7Pu2Vx9jaeIyNAcW51GhU0U9XKvrrMyXexQVnOGrCVttIsb
uuw8ZzYs8xyC8fRiJXrlfnUNaFw3+cf+88MC5HbIKxsnYFjJN7U4EulyqtDsnehw4Fou2Tmv26uF
NWBKJsOJMTk4Gnjidf4Kie+DgdsJHCNk+3zhGQ7lTBSY2MT8qEZVXUltlqw0GxaAnEJYU7cDEZex
1JqHf1gG/OlZmHZn5QtN03Sv63/AkXDR6JcqTqxxv8aFqxYFM8ju5p7lrroJpEChxOK7t8Ow8EFC
icfEAkuJCxTRdLLdjT90avrcbzcUmkXRmbEZF6JQmlPWR2YWhCO1nljecenQqjIwY/pCOuh5GiZ7
tR+dAyLB1UaYr8eXdyD8q/2u4bA4fyeb/vxjU/yo96XT2O5R9YrRA7t+Qi/J9i5Q3nbAUNSKEn1Q
r5NOoctLU+nIl7pK/+AmU3irRTzXPbQJOg6LkmveoePuSzChxoO0nJ2zr+qm75sihX6Rpwj/DwbW
g6s+9+eFl32izIMZWP/Txib7WrWzVDkhnOg3U9BTyir/WG6qk22QrLy4vveygDGvO/kuKtS74cl4
ohG7XRvPCJcEU3pxRtKjohdlosrsMVulPhXPCgrhHJ8tiJ8iOTiaNvUvkwBSaQ+j0Mv73s14HQvj
dBuQTueNkbAyNGPujisTI9N9beQaOr1ZL6pluywXcliIsDg9Voz8jTu6TPOhV13XO41/zu9P4kMA
p7sGsVfGTasWZ2v/BaO78O52hqOO5XraF9bPo+gq7mcU1m640oSmE6YYD2BIlaQon6jEUbSElPUA
uOwkNMQxpktDvCh4uGl1+upoq+vPehUpLbTy0IRP9QJfCRFOltEmac0AEV+fw66NdCX4SVichxAD
p7Dv33RnvYKgQ4OwLk7DX76mvXrmfZk9SSZVouRHAj7bvaFi4ZtFkNK2L8yZHL9vzKvpPCDlbybk
zir8cL4CuiZcYwI9+eIBkWjY19cR6lzTSSKn/0+6N18XN6dFk3EUsQ9UTdWClAh9Isx5GjnH2lrD
qayo/5bOh7mvY9c2NkcdqvKSK8p3H4E1HtCJ7ioSCVX1Sp3xWxhciF678VRxFeKBK8SM0E/67jq6
cOBm0rwSVK3q4LBrJ0UgOQPvvs/ltBYmig6cZMpCB0yWnI60K27gTDVRwQxVtSBR+zC3yVn1ONmz
SeI1RvZDhTHtwy1A+QlVj1gfY9ci1RvrhtMT2b4eKJ4U2CNQt4o6sNgSnGqWo6xE6DYfFSopRaRd
z/zy3djWdWhC/b/Nxmes4iLoYJ6AWNB6PcLpTJijfkMSiGBBzDB/8cfCE85ck8QDsD3qzoxl9f+/
uPtyfxJWMMD2lLHlA+c0Czz4o3ZRG1SWm0Z9nUEtHw6LAmt9wAzD0HhrmMewB8+hy4mK6wEPdTnq
HAmVNZRP6B26eghmD8gPp21rAcWqnlMPmmpvuwv7M3KKpWJbn8rQC/8ORmSmRa06AhThWbi/slk9
xRdeuFsdko85wDDqelwncWxPfBLNGZG8MwwpJqylrTcbS5AQrmK5M97N5siAz7TUwpIeujRGFCST
mk+Hts4a6a9+S/NJyXEigJhzKf18nck9j6XP2Hm5Pc6NU9dVSViUXGmxVsmQGhTu0DCGM5xaAvXK
yffobRw3cM6lW60gybpCqi21SEbehShsBuh+++8UCeqd/GbPYpU6cFO3HJvqYPX/Ng0dodYJX72g
+2010hWBN8RQf/SZyHLhPG8f3dbZoNcYPa9gQTxWQLSbl4xfpRKSEe35ds/tuds3bxoD/gyPtv5z
KMr0LYjnhQ/J5cq0GP8lGM6w/YgxkaSnWzqIFdeaGqqbcWpgY5yJaQ3xDo4VwklZQ06f2MixIKFg
yH5T5VzhKUt91aLl6+fQ6WqTQCViM7bHgR+88QormmNWIHeaYAY51+QEri0yk/vBp9AtiZ3xcxS4
3Z6CvnmQTMcNWD5wv658OYyfzJ+YHeCsGBdH2w9oy18huHZNqC2eRfyFZWCLi0Jt4EwTxye9RoBz
hBR4RD4nOwy66wLhH1d/U2z3Di4JM/H8XMiQtSnCOks7Dn0rP5hZjO5Ad8NQlvhiL5jM16mzeyYx
0JTWUO2yzSZ21r8oH07lhKCoKaAwrGuWliYAmCx7w3Wk04+3uvqu0wBDhDSclxIEimDSxNnYEqeb
IGgqVIqI/32hUyOPUCdtjAfjZOjYxyHrC4B3rd4CdHWhDmOLosxz3znIuNHL79R0+ku5yFPzrBS/
j/zGGYEpYDubmN4NqvMFaZUG3Hdl8hU6CZmzr1MaZom75Ucpq3DaMGZxRQigecGuZxwv6+O8IcXQ
eRHBaWTTwGDJ+vM1txTDWzSXJAzYGCu8jubpu+Z3EOC4ULUpkqmhnQi7c+77KLGFgly5jnbjf6PH
oSy0nSHXvpFjWSxNFmnw4nfSotTg7f9TknvcUzAmUvPzQXVu6B/anEuRRAKZhYLFSjD3Iri8KifK
/g7M9OIlBCV/GM+XISvBHFlM/IScB3SUKWqWdpAxehgxoO3r+yn4LRWy5FgWMulRsxqnnahscwa6
BpTy7DcmgL1KJq4AO12aRBIy0gqlKhg6qQwp1FBZoINhYbNvyURJV56XJahwrZto/wp3522lDCvv
BTH5lYEvYirhLXp+2mZU6xiFiGlRgtkx5/Ss2IeoZ1YRhiKEkhPyD3GgY13IxzYyaQUuCc987KhU
u70GTIQEDGV7337WU8WU2UI4GUc+dYeDP45e8ca+zzE27o1nm7hkG91ZO6O6Nm1h9OwY2jiPxgVF
ZunkdgcnoEg/zglXVdsvgiVrh+DC4QSOQ7C4oxFu3t9W1TmEll3w4PYAm1SyT0cil9siKnd4eksh
Ifc9rcj37npXjWa96/o0L0VzDyqk2wnHxiuK0LOoleNJn1g0IahhkR0bLhAJdzsMlfWBfqTrRSVn
BDGo0qw9WANKw+vY/K+gwldqotyOLQ7XFo8DsZqTOqY4mw5tcytCJw+oLbcMSzBxzBECdofG2+QY
UrjV1CFP7ruMmBTfh9T9ITHB6PL3YndYN3AdQpr29nRDX9jDm3tY23Po8LExcR33FhEjyFhJmJxU
7TPHFGJBPAE3OpplotT8uSlb+RMxlShlvdSrOvaeV7Gk7N6U8YWxUKxv/poH520z47Exy63OcY/Q
D4q/DeYmaACekmKqHDF1Ar6URBhbb9tF65IvLcCQxu3qb2uWHh8Hitoyx8Ibp3KngdzLxK7cdw6R
D4z/Qrei60R3EMRw+l69GIoMean7wnTAEf7kkJrIUnFQKARDf29G50ihbI9lMyV/DL2jasFVQyMz
Pr0+ujLx53vGkYLegn3RC5CDanwwFFfCuOif7L3vXX6rP8h2B3is4iNenBRlvwC+T6B64etlwKvE
F9TMoli3SpACtn7L/u644R4ySucdMYWAwARj2A+1MptprMu0y/3GEtZXuGyPy4L42bdViA1FUSVx
1KjKkbevpASSPim1pMK/xqwkvT0h7b+Qff4NqVKTJKqhpb818rOR3W+YMyt0MB6j9zfWgUV+Yonk
vxIg7APQ4wKDtez+92rN0r9sXaw+jvKhl7AaClqsR3ZjkT3dotaSYYDFew7sJN5Wh+UOY/jTUlW7
QqUeF1CNk68sOFOQ/54pAQ2q+0dB/xBdUQX1MgZv07ZkUWHgYqa+aVOaXBh0G7hzarg/W0lwEAfe
JQaKrWxmmygfbupvon/6e1OOWp2f4NeLNMcwyYx4IGlQw7XFDQVXF2hBflXMqt6x1MDBQYu1odFE
a0NclPLhGelopQCi/NRL0ppKz/TE1Ci6tLB6emJlpyqFbrbBufEmZOw7UuxYWfj75pcd8ln3qHdi
VY4xPfL/0sFAAdKw8PccRKXdRC6w/00+PUAjOIQTY7JmEnilaumLJgoJhMn0AJAZGJi4gNpNil0d
CFP7xt3QkNNiRjaPdjfwl+D2JY+hsystcfBu6F6QFO5fr69d6rWA+FLqRYW6yd1DiPhpn4bhnXfx
o+JDN3EdZVD6YpFmkgWSIQebm7xziNMYiq6p4csESGcgXuK3LTayPAKkE0v59xDfoi85YSUAGxeO
LNZ6EwA1RcbxO4UHiLMIXlyfRpVa6p6LHZ4IFMs7eXB8cUj6jOBq+n26+S1V7/Tafa4XONJK5GT9
6gkD/ZTYJ+fn8w==
`protect end_protected
