-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0Myv7tyU0nmIlVH1EyD01lUP4TskaVSYhRtIrFwEZIgejdoitlaQLTwC7+Soa5FRLbA0wffabqZN
BDkExzAS4RCmN4yn3g6WMm+/T6wEHvRumaVtPBZKRC+yqLF/anMTMuFo82U90iYwGC4iV8rWkOx9
ubrPRzb621LcE00TqTs0qtmaqJICxsmgWx1DmhrzVJfBdWG0EpiL/TefGK3zH0YWTMfCD0+IETLj
BuODRsmWiKYyh4lRH/kthjfTA5HZYQJTF5WBafOrPWDqq0UC1pf/61YIJ9BWBtY+Vdg/vZVFK5SP
9Xb64MtzIKm85NSmDPu2XP8ayZqM6C3K3/k7hA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
7Y7RvaNBo72VB06tc06H+JGjqllxzhNFVpSJNa11uGren6XJLllEZ2jTXSGDl5+AkmUVMdAVVR3Q
N3wFP4E/bhZ6VTuiRm7ncYaDXI+fY7Ear9/qlboxjDoj1pF5gNbWkvBwDDPgOIxFuxMhfDucsmLY
dxr+AkBme/d/81ZA6O8KcOP3YyJetqEGKxnT8q3G3Vmx7xIHKl6e9FcHnpkljGCIBuUGBBHhDWvj
s16BnkTq1CbxbedASKEjpyaCUIaXzz7M43wshu4MuORA1njxm39V8iuh6tsNVqthpiciZKd7Kx+O
vArRZJIgbB3pUtyFQV2Xxzbl4ZLQMMtdDIiOyh+3Jw/50wb/JJctERqfsyglBTozYzBvvE0X7odh
XZk8ePJ5ol5sIkycFLkOFCohUe3R7TmEK2RnrcRbNbTvL7ZNB4VCjiyTUuoWfM6v8+0slQQuFdEk
maOMcsblfkgVqOS9e9a3In7JhyIGJ1abama56LzS1bMJ7u6CHCZm4iE0jdfK4yCsucoNZ3Qsc7Fm
bv6IIrW5Mkk0WgokaZQWRwywZCgdPKTwIi5gYAq/c0POxbvUkY2pdS51fJ6OnLEhol1EKZuGcYJ4
pcKWz1lUYvXhFAxKuRAi6ssFh/9S4WS78XQom3EdyFAb57Ir6ezwgiPOcAHp0FT/8GqfewN81yP+
bcqbI+lcN+kHXrC431htK4B/cMTmobmKSH1pNcAusLGK5VUzykPasTcHq+0CsMD81xHn0/PdZkAW
BsEgY+mGH6wMWckrGIZohESwXOTsLxcN2eVGphZx4/Kd4Bcr3maBPrM/WwjskKJ+WRzTjG9d519q
Tr0Af+9lHzjIXLtDemxSvn0Ui7lMC8Jck3yRui9XGxL5xACq2UZJwkpKZgRjWgpk9gvfMR1B+2PP
mgh0XTQBpmRnpUhRHMCKK/wkRgWLR/Ysjo7j+XkSgiKJ7119YCDcDdRLWlK+sk1O1iPJ86VaTrdi
RZ3tYr9UtkBo/kb/xSaU6Uo6QuBY5cpgQuWT9GsZKTbeW2Q28IVD9Jxdz5bGcsyd+iM70D7SMycx
Ivj6CQvLMxKBlAEWrav4sGA2U2m+sDmIlfdcIhUfoEvsaeqXd9XLei3eSxSoVLoWBcyxLInR+RS/
+8X81dhMvNJVaPS8GDw4rcGQLXEMrhAQxgX0eAhzqN1hOALzglkLzDj1k80B5bQy5TsGB4STv8NH
BTT3xyrs2qSvr97tIoKdo0ZXX/+csbWOpjQubR3oSLUT4MvlRTx1ebMfp1j9mnIHVEBmBuimk2Wt
6XnY8axh2gu5WTbGdMhECUW6xseObry8Hw0HcGZjSyImFaiYYtF2RIgbq8tTSnwKYuj/U8m+RCjZ
Vzn5N44av7fWA5NwUMew7+wXchBBg47pAdswL8YlTahMn3RFRXLK7/uqty1BgoT7hwkS3QA5Ya49
gyeBa/j3dAJV0fdkUvyaqfg+7QcpvJJwJLmYP4lRHCkJ8yGv9WxiqIMsT0V4NR09MU4yNYp/tsPk
w+6i5f1VzMb0uDEPxYSU5/U7vtOkR3elcD520v9DFTxpx7hYg+EwTkMFSuZEa8Q6NUZqlesdjp1f
kKWo242coQ3+9o5g0ibg6A29NCqp4sD17pAVl7MA1v/eZ7A5nODoRYJRkS1mX2G+QJdtA8mpmS9H
s3Chywg8xd7kl/uV50v8gm0o0A2OlVzUconi6JjJ6zFHCFPw7+pjsSMEz9Zramqeqnw59xkvS7/q
5mDOLpyKBESF+QX1Z/G/GXkrQ3daVE4GJoH/eGrMmXCSegtTOg9t85j+r4WKtM9qtVEcn7jzgAMu
JA8E83p70Y/avU18g7LkD/ieWzg7N8zllRYYFAry0/7FCKMbKH+ideQTJA2sk4cAyhKJRC3LC9s6
9pwJzpUOQUqcgTM1bv668qb/pTKfbhEZuXBtpVeOlAPZnYHsUg9HNZeVys2jQ1RBD/6yldq7eOGm
U1MGnhUQSvBJDs+z06dZ6e+T+z/XIJDyZ1ReJbDyNCYgW3IpvNKx+U2961+GPtz+oetXGLjMNogX
99Q/V+KMGM+hX/MDvQk0Mgq224tBdq6JKJ3apnVpbLLiICgm5X6bvolU2NwiTykK3Qu1S/Q5LNB+
JEw2k6d2qH08SrUxhcfK1cdMsYUiKyXwwkGdH5QcC3mJZzMyI/QFShk/ImsecqO7WNAQ3YRGlh0G
denA5eaJon+o7rwXQIjovkxuLY2uQpSsWgV30jIfqWe+S9KAdKpTBu253FrB8QATiyVtPZxg0Olm
74XcimXNcLJ/aDn7iYpsWU9hNsUqcuh9AFBiOcBew5Ikzep3GkBKOKoIXx2jlN42NOb51vKfeQXh
wMabhf8j1TZO6rBeE6qvOR2V81VhNiivAEHY2i7ToYlqc8XE178CU8pTgBRztW7EL+pVqIZw6Mza
dp1wUPyM7Ios9BUBLty5fV4djkraBCpXTONuk3wcixCP3cal1VOYOeXHF2LhUYd5EMllfW6CBqpJ
rmD+FB1JoUEtZKw4iwnpgG0O5WjRbe0CaB8SC8XfGsDFKgfG7myBuBRiE54NKsrMbZ5rBQAec06G
f218xLjh9YTwmKNPDCwWBdHdeztaZNd/xefpldDdRdTLnw2Z2UD24lCTfEKyWogvEmziLYWokXB1
PuPk9MSh97Ag906TgK+bDJ2D9Qi4oCHRlVXa8Lb7gvSN3TGEiuQykBq04m3Afn6EDTR9Ei72/P2M
cga1IvN4WWmIttHXHPxdemPID9WBMb/EMuxkfmW/jRiR9oOi+6hWbs7kOEKO601nIs/hTZgAHAt/
8y5PW0ow+o2YvMBJ/C2WnQce6YVy4X+ASLp3b/um0B7R0bMWMMDAtQjabos/v0KBKF6KLm9zbIQ9
s2+CuV8ysDziVAoVwxHGtoenk7goQ9aTt8NevIrKxhqCIApRDCjbGwU+faIRwkxSMzUOg4BlQsrg
5Qb6KkjQ6QhxrK39FeQYdb0Td3ulXpWSRcRR43TE60DRg0xQQ0of1C/9O4dZRvX0sdMvlqYX8jP5
/wNqSWcW5C5iNSSI018KZ4chpSq2sdJepcXMGtkbaGprwGNsXmD7PVRGRF5p/17bC5d20xHLD1wg
Upb+dK5kwsYuDlAwi6As8ByuNAMRxkuosSOZXvZ/CDsQURzjBrVvhqVXJRjy9MZUx8LqZSA1E2ni
+Yx1rQs9Q2K15gkLvByV2IEM37MHn3HL196xK6nM0We4vdqevQEtLCOW7Mia7CYwV5aE87gJ5Zbg
iCepPStEqfbkeC1OlgkFRhrm6pDdcqGVN/Dprt4cqQhf54q258eLn9gIFbsnL63dwgvV1PZmk9B/
Yw2xOhaEDhD5C5ounXuZJ+ycH0CB3RtpPFhJJY4czlv46pLouToiSkvr5ESnzXkmR7SViTf4niIJ
dz9hq8Uw/9mWRRTG7mtq5v+5l7E5Tmd0RMh2uqEvuo1TfRdzmtqNv+LnalwcJeSBB/lIkXGmfoYd
mN++0Q3R3HMhpYTcAySdJeTiTGnM+RzycmfwYoHz8IZiDewYBvjvcbHJH/Ix9zTSiaonaiMxm3w1
1A5VyEXq53fAYLTYfY2D81xU+tzt/ZTjUyoE7z93EBUmbDVeptPPc1SnsNce5NjtUHPCcQactsSf
UhSXA43DvIbfKRKDVZbL/J/0+MSXYAKpb8jySsDm69xw3k4kxtxA2Wu2as9cOyGuurCNoS4dvTkp
4w3F5QwLod7FNHK7pkTUfJug2niztZXKe0yoteoURVH3rBldX1os+4X52hqAPgCT5eGxz2PqTtG5
NVARLowuU7ReFu3kVXDoeVANsn4g7AXXImhCCsGnbiKKTBQs5Rw5jcJepZF4B1U5QVPDFMeIrW2/
JK/mrfXoQCsAq9yq0lJJ33kWnFCpwNzgT9ss6WmRb5rWblk1qrOPcmQaBe9p4A/LYR0kbtTMQ93g
2EWFltRL/VM4OI2uuj6tIgkOcG3mExRnMnNB1TjxQHf0Z9vfxlVzT2pYq7BlYESaZ5W9Xa+gAibs
oqYGYjcd/M0j6zEJHLoG/PTdi8wiPb2FYOooJd+ogI1fpmSwGW4KQQQDVotNVIcGvPspz2jWl2yK
VgOtgnqGXDE1HO7nNrAZ23x9GzqrNWowd9+Ms65QirNkzF3xH+7AdXpatkq+6V7eDsOedzQVJgnv
gjw07IautBvhoNszdFvPcm855k3RdEN8r0PEzLZj1pmdgHr/1IXgfBN5dxkEXci88rjcusWF6vgr
k9z1xlbu5Ewr3b00gNDZCPEq+IbrXmrqMrVdb0w4y+jffCHiCzyj8yInDpDap/QS0d37fJbebHxX
7uvSt3pvMQzv4Dm2FGiAbzegFV0so1rsG1d0rxk3mEBF8XSGCe0K9esScL0FY6m77W594wdlTgnS
zzt00XQJ8qVt3JfAjtXpGReFURxc5A9HDs97K3J20KjgPOCbGK3jFt+pTHAtS2jNpeauuqB4a2id
2JzByrM9NJjkNtsTfwECcH5yAUL8K5rK4MRIAFuDLkydkCw1hyrkBEhsG9naZCckCd+NkaMcX3h/
tc8UbVFudRTPlDiFUZ1wqJ1VeSJ1oFqXsy6ukz0MfTd/FdTG7BI6TnUXc5VvyEEXq8nZTPR3uml6
J1a0G3dF50MOpULlpsVqwBvAjMAlpWNCbu7qStyobdorp/sOUCaUxLkJT4c+hBAScHQgW20Pfqa7
b1f+jhxiEAtA1DaCZuEb68toZ7LgKkicmm2PKsemqWyZ863dMHASYKWigx+2NgzC/kVOc+74yJDr
Psh9/qguUIlHuqvz05txba71KG5N9KoNxdSdWTgGWOR3Zc1cRK+awPIkZHV8kaTfPTwqK3H0t2UU
xtQ5UD7Yx4i+DzoPDucIHcINDp3rzF3PhnJ0E3aWX5gIaKa4kQI7Gy5E1iRSN12ASLgbjmsmFE8H
+B5PdIfnHEjQsbpF9e8tBoqE3U+419GHNoZoCuib98ibdaxRacRIrMpB73qxiZnkr4zY89oE9hWN
dRl17MWMcb6UnNaD3D0QrlrY5ZJYTLyh4JnFDTe7BPThrhU09h0BOew+/ABMUMNKvjKyayK9ErzW
fbXC125BZa8HquWA7cLQ/FkbBFgwm02+Xv3JFOGGq6dclUN1euIFym8Pm8Z8FvjYajOw2XPH3iIa
+gtVcMvU5QqhqhBEE/yTB8yUKpV2fYK6kIUIsv5jjKlTU8ShTwLCPpkvb/aNhmtkyv7XlfC7GwVU
x4U22kubr46UHIF1eGu0rbYqM+nbY3trxjhLJMu0x0uYn+CLU11JsbuN0bEXjRgWjJpMfh7pGheV
bL49W/7QrWI31GX5FxFoD1aezeFSmX81z9vBsRPmZwZgkcofs9hKElZ9lf8A/CDCc2IHhDXzSWjb
XjQGvuEiUn3bT3OpHwDgGPzdHkUJf4hXJ+HB2sm04smDXTIYkBV8iIfvos+83vnoLmvEEepp+Bz3
yVFIskt4xsi6VPcB9B47UTMPO6obMpkV9Y6CkUobLo9vdWI9YVwlHkr4G/OE6jO1vetxtLzjbqOq
Krb+T4lKrkYDfAttCC9j8IS0HQ0G5hTKuVwLS/GjV0aJXiKIujBnxVVCxi1BZ4TLuFGGhBnAWqCq
mzW8RnOex+2P6iJrTvAqk4A/R47Fk/beEr8PxSqPbOcKyWH6o8grdUPA3n1Tq2PKBITjTv6eU5VP
ggPZNtuXkeHhah0ZlTLqXqz8fZl4/sv36H75QJGyQZTYsZyexfwQ+NNLgcLrvmtQ8gfnm6NZ/YHF
Q6xaYPAo844YLDpSvyzRYay30qsGjLl+o1E2xbJ4OaxJeZ05ovNTeugko82GyySdEq9uJ2y57FQm
tYy6wFJW4lORgFF1zJ4udrEdNncEVw/Pn4IuvLbiuM6ep+BUAE3ITcAlACXhbCMJIN39CmuuL8yd
XYpmtd+hZ80tAlubt4C9VAYku+FD3oamekxCNyv5NU/yucviux+5yemOaTtTJvlSROPBOJMeQpRG
/8fcXcjtVQNz7p4/7qYAYJH/8zdmk0B4Uxnkeg3T6GvJiZxh9LbzSYlD6zL/KDbWQchHOjOIRAJW
YOplAuBnHQcdvdu4DcYjnOmFlAk8iFmmJGLBzDn2uSgeAXQly/biR0whUVLKUTAT5t4BaE1vmirS
FE1QRTINjcRJSKdk1UUpFX0468sxRnckRQXoGeSMzSSG7TCZWIVbs4ju7q6wI7ue/EDTgRwdJz+f
krHVzkfUt3QnieptMg6yq9+Y8ZBtW1Iex/8JTruG3k8daN0b2EtfzpAPjopN2Rg3naNZ4D7P0+Kx
xuxOHkBriOmPQulEPrrUSKTEwQ+DY6cYW2sMm+tPyyujGaTtFgSRlWcANtEanPpjI/rr59J9uLlK
0d80MQFHCWjzwknDD6tlsIp0mjl59lIhAcdf/kF41aLIRLDnSeriK6S+jSCsKbp38PYTHjR4reuK
gHG5WGP7xr+AnaxU5xnAaYmgnQjZy4HPHYTuQMhzsa7mCNlSGMBI2QYzGJ9QLYrzvHV9umJtMy73
qISIYk6XHIEMqfxuFDZIhHXA4ZNNiB6qMfHOn+1k/EYmczg8SNylUj4gy1HA14B5ahgmZc8z9C/m
QiR2ioO623EmeqQKIbk98wDzfwbPSMnp3zTVOeXaCitROPNgeEjElsQvhuRPd0AVJFmf/BWJ0b09
Yif4HcbOfs9+EMU0P/0vjiqLePjuH/KxdWBig9F87PF8vMpVNxgXhMvzdurq7QpuQEreuh9krFQ2
KvnVdgVUkQZc74lzOXdYOuTxH8xv1yfn/Dk0YGJ73yW5588FxzGQWZPOQ7NWrOjX+CL2SMU+renJ
cjb4AHzQxbc8YZQuW6bMOJRD4rkaWA/i28kRGQxArdc25WhB6m6nU10QOuiLyUkl3mUtmz6Gz2+w
CQfFyna0fUbnfSf4Ch/EPu9w3oxLC0w5qXLOm01it9yHA+pOcK+41vhRhaHc5FecAyuGlmYPVMbi
DgqDbd2YexcO0WNTc9d98drB2zwPa4NMASKwqQOf5CyBTQZXeLCUGNzOq9J5wMeCG0K1Xq/uCxR5
b2ILTKx2GqMAg+Zq4t5PnZBugLRVKyr6rjYXU4n6/CGQ+w2MT4kc5qnhlOfnNRDHbVcCmtNr6Ha7
z4/TcRub0bK/ChtvWUBcVTLwlHNLf1LP35FMCGxeGkfxTtCgh7JhND8amt66ITrknFg/cgX9nS0A
Og5s5yRo0rkfj2CHz8F6+nJ6alGHS1kEqQ1ARsn5d7/7Byfx7xT8CD3cAwou1dqtRr6dkx5JD3kT
T27YmerN1tCikL2HGkPN+Mleq5UYow5Q0B8H6Q1J/n4+SWRHICHFlgjzczktEZwScaCkUjNQ0RPw
sCcBxLK8uT6rmkT17j6sR91wmvFk9rGfGWS3TijcoZ0zXJ9raWWnqHM0GS7zi4xW4BW8guFKesc9
ZMiVg019KwWX+gyAkK1/nzJwzJDZHPpEMrwKfeyCLX8r0HoGe7XtktkLo5vwJ3tJhqZijAo3zcQY
LQNxMj7TZLJcS69g2SEHIIdzebGRX37Eg1eSSjSYryqLlk8T7Ce/uLmSFXMphqU+UrJMI0HoZRJq
NQR7nzFOS7KBrPnACszaf1vIkFgel6J/f1Xpk+a7n6IMKvx/tLr1KyWInpLIWNERM9UIAeBY4ot/
q8TtVWQ1+rTOyRTZLL8Cu1Jc0UubwXbddM8clBnkdNRqMnyvVd3ZmS06IVeXzpmsAO0H/M97pBWP
XNXS4mPmZyxlX01TanWoKd05W2/FyrEHclHVRsvfjElTZtwVL7r8qowbBkef4TUjffh33x9oRXyT
xF4Op4I3ZIwM1ApzQbN9HR0BP0O0kZNaAhuWgwweBcAFkCY3gOOsryFTEAA/wGQfF07x9WyVZX9T
Mf/JCm3vJz2198B9cmdK04rdJIT8BUktkbciv4KObwx3eUM7gQcLReLbRiOEt5GLT/3BUtLm9bI7
B73dKNl9wRwzOd75VTVyb3mrLV0mgAYZe8jyb7xLbIpqVJ8mKzzwB+XEfbwoQFRSsFaJQaxAy2t2
8eUpQBNyskUMa/ZQ4bk9JcFAO5KIYHdyODanhGAom2+jKWkMtwIj5f2crz9Fw20DUK51tvPKwQXB
qEDUUtMTlN523di1UHPl0AbiFTmEaChYgnmZh4ncIT0gLu74aS9BUc+N4RPqv8NmOBLv+Lrkc/Rt
gmdn4XucTPjlogXMDun4syL071AjQbUlBTMnuh2b1Se9Saa4HgaINgwY+yPLpfEjyUf/h/8Vn74z
VWfWt8UMARBf0gVxYpVyJfd8UhHbAV/pqGIV01OF4IskGs7K+I8wV+oQfqqhoV+TwtFAYs+ZX8u/
82hfPpWcoQx6RmyHJmJOwcfJ2Y7RsfU6OirA3UpEhx0WAMzYojey+g4BofaRb1vBqll79mWkwBFt
8xFDjTfUuhiho92zXG0BQ1KlzYzDWz/H9kvl3svsJNuY+IOEWLXqVghB4qESKES2cJrX6R5aAmOM
dDV+Y97eWeKA430XuRFN/rRDPhzxQlYXC8gZlb0TBTwuOAPpsgsao3eXuf/YENcxBv8y7OhiOkfi
7mXScCTJM7wuMTFUDTJO2t6SdRYFwvGgJpx6jMeIXSEofvgqGdJ23YzBgoDqWwnnl/u0aiIIP6vZ
u3sEBPXF/ZDCF+IwnZZerEZWDrPDAxwNwONiNyxmxg32u4jsUzJFboBF+pMTUlc2/ooJVT5KwYFD
BcjrHoQjaO6GgBrPIqCCkz94q1S1MZeWd9fSVtfLSFHebbsYbfnvuHSeP0WHIY6PE9zr/EbbJ4cP
M5xuCaaY8Vp3w1tBpEXPEucqwZWq9t+ELDOaeRgdAX7wawuvuZfDWjLRFD+al6nC99/OJYyvoARq
ZBfJ9x6P78Dnu/lxW8QrpIgDtGWs42n4Sxhleqm9hKUvKmO4f0x2U7os/jlc35wAmda0OAoXGMxy
JJI8ebBmj85Cn/cTdK0EHzlDO+srwx9Hj0kZjcSrL6zgU7+BDwKpbU6rTxYCbI3rC3SF2Nsmvvcy
iQHI4MepcbmMYXl4eadevwztmPx+3l0PWhPnL5Hsj1xCSycMjTBmf8QYnJwoaFLL2JL+xDgq4t/k
y2FpOuRyzB1ioqas7qhayYJ2YqV7MjRHjIQnCmbrD8KPcqI2MQekeo8z8m6d8DppNKz5pDZewdIN
f4SyAz7DYapR6r+/Y6JTnZyrSpkIq1X5OfRhLoANk6CEZJ5pmwKdT+iMS6j42oGle21O9WVl6/Bd
5Pvio20mFUuRXMY1Y0Fol5t1zrz0pc7tt69+1TlTOrMvpFENbd6VZVUAQK6VjZsL+XWLWOxdqAEx
x7JmR33VR4SMISeb43TA6XGU+9tVhAwKXoS5yiVNpZKsZcdzmPlqMKB262FN6vNxwlDkl5dEzi8o
NUSfNBC+zIjhXr75n/ynyZ35mH4ZRU6ZxWQJy30XrqChjiPmQLtKRJBPtmv+IkbkO/cKNrxJZf8c
7+DIAHxdlIgfsGUqrvy9EFkBZ/hNaQhue6NL4tA1gft/PjrOEYM5av3x6fTv7P53P8gJvqe6oDpO
UoDSNTDBwgf2QLv5ECEQ+yo0ZObyfAnBLDYxn4nLgaShXYM3XpjOhwRgahfv2nPqhQJd8Jt340Pf
fZBSq/q7E57ynUoKsw1TgPpGoCCIlm1BN+/Rz9fcTSkGRVDuNtdEbtrMFbdOsAAkHlVEQN4uo75c
2VHKNo7Ufn5qIBVRRHRJpklk9RBt/BfP7YmidEtz858RbvuDpgV4rBplmZ3uLJ/V6fh+mm5EWtxy
B0BCvqN+4wziGQ/hNXjHGj6hBPm4awmWYjbvinaGEvdFArDQgqYaSLAv9SNjJUnP07ADnrXYjKcY
6ATvVfDgEaX3fmAaDFnNXv685QrWqR/KD+G7h8Fn6Ws1dic8XJGzrFOcVD12tAihlyjd4t8xXmJa
doJF0tYeBTk2yf7jGw3C2oPhj/8EXlEPwUE7Z7B85NJmYYuTwTTErIAAfL7WbZ6aQu+4q44fB7OU
6KGIRuEdfBiM0QOX6u1fXf/UBZDQQmsud7UlJGx2Y7t5jS5QMinvol88rQ+Ttqdrq8Z8ShzHDtvX
Vm463cmBOGcJN19ET3Fi9eyObK+exXm35PkXTcmNAI51MZNCTy7GUI9lbRFZp53C3svfAj3Vjd3r
U2iM9Bmib38PXR0Mtwq1ThGUKXIzmoLxqUuyvk94GVrYN2ER2n4uvg5M+Ok6AS4mmP3o9zOEf/Vz
DQ==
`protect end_protected
