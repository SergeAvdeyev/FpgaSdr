// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
E8Yq5Utm8VdsBEopG/nJjeIQ0D6kyKPxA+hWTmXgIzt0884QW86uTkypF41AvCLhZTofXcc0gFot
0NM+G+eIUS5QvKwa7yThz9SMTJGAN6f2x+9jmCapGyJlUzHlyK8UtXkTtiICOYCq7QAWEwKVC5YD
qfpfe9SHEVB5s7ZBy/vSI8OgipvCHJN3bPRKCO1+WcLicM582ULm457z7IdDJQy9BixfCpV186Vi
YN02zkmNBFVmDKx7i4nosZWTK16pfMwr3gjUC+euM6D3LOhezRv+ITeKL0UnfR69Vb1TvgrN2zPx
kMFf9fTQru6iQuy+i0oC57RNu/vGZfLSdJR98A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
6elZV5IHAWT+k1DeNLYakgFXKpeeTOwtiqQLTEzn36Dwe968D5DTwNZR6UvBGTuZ9gUZ4ocngucE
sn+F034DZpSbwkPa4tKt3fSSaYDD1I2iZ9pUCjKW5H0ZPBeVcVHkVjUFk6Nt+W5KJfh2AyOuSMPz
Ub9BdXqFOUjarS738KIyvvKmuqpDCUw4R9Oww5MtT0gffTilngfheVJ5HlRaZv9PQXAWnF6RTUiP
s1eUaIcUCTHh5i9YDlo9Y7OXjIQCPLqIxXutXFxTu8cOo+8j+/puIJ8xbROfHRmZymu+hpaKB/sc
zHphZZk4TcMilFckmW+1KsHA+co8l7LvFpsr4GrrJcXEe2H8eMaNFGOpHe6bXAHjTzwlVIsP/ztM
a9ktxL07VUmlEdD1uY1cIOM32LQELcee+09J3oP9IJFRAtuc1beCf8BKki5NX/BAauchP55At1Bs
1VyI3HJZRogXe0y8cLUGBcYqkc8/P9NTA11c5eZ3N9D5bXEGm4zETbBqZQVt9daJfqdN8zATZs+8
zDc9Usl5lldGcPokdvU4l8aaFyuQGhA+9YAYVZSMU2aWQG886xskMNjN093i8ZMPM4rmiIoWyFU4
15WJQRxvEGy4iCBdOGEAHyqBNxlcsTsFjEDf7FnVBRiacXSfCmCxkCMRFWqQKQqGAp6lG+zkTFnf
6ejb0haVSi/EWkqkRUKbsuPqnJRvwMNb0x1/pmHiyU0dkhKcMis2Q2sKyMtRTOvVu6hVEfAgoUyD
mE/NGVrmn61bUBE4Afp4ivQ/o4+Fu9y6hFHuY4PRUlARh03zsa/keEB9U2WQWkm709t88N/SzVVi
GUfWkXRTyFcr3PmdHmdlLMNd7u/2h9pT6z8pfvVEwZ7ajShNMH1p9mvsXAyFCWCYgdHkSV9qjBGr
aamnKm7E66jzJ60Z889Tk1sm2yf03pAlSPD5Oo+xC4PG1bZXMwCXP+cjcsz2qfJjebM6RXDh9xEe
bVHJMhaK2e8AwFJKrDSo/xmvWhi6nH+wlfV1eMvTLOfWluTxARCT4mhJroedYQOk2qg5G9/BF60s
ct/DOzVbXIRF4MiFkjnvkrrU9weGXwKKZ88zPNQyT+b1WLIMjk1Gr5u4tWaktJmQqI1qp00v9hV5
VUylL8kjeIyTdbyRMysSprxycezkrM3OAvsSZWsxdJPREyzyhXW7m0bSA/00Fm2ST7S36ZvNolvG
VMqOry2H+0DtZzDdySrKLrePN+aX7xc2S/v0fIlAxNbF2wkZlCv3Fi7GeBCN92m9dH6dLDoLE2ex
Zf1LXJXulKwZvDGHrjkhBocSBPeskptfVADYB/1yyir5hm+y3CdyQZPmFWlYrhH68sUyw5iVwwPA
GVJhDgtzku7Tm13+LdpWggaDC/SGuIa6RY7NKlRnk/Q3iJQujoKlurIeGmLjRYijC1armPHv3OiV
KrG1DRPvEqx6LIF5LaX7r+ja84knqP0bpSmjq6KnzpDUksD8wWZl1gHhXknM7pA/rGQ+piH9ZxGS
+s38G1nJ5GhTza25AuJC1RaaAln6sc3TdjjybrkCx4V/4N3ISDD7p41AmGAeoPZDh3qEExaFylZ+
gfF/iPl5chEvOppaDXUB3iOza+KfSo7A54otv3w7c1r+xNFKZkooXrk/46awi21QAro2gWe7/Xry
0CC4iQsC/9LDAeiNw/grt4cZH/lHij2pDPSonsBJB9BXxU0A0/iPGdSybV82i1aIdiPv3SD68Zii
tGXfkoBqe1w1awFWqlZm+GJDdBIX6hqyzh1kXtrLFIDi3eLhIA2uhiVjSZICYSh797S0E93cPJ+I
SwWd6325CsAp9I497wjJP/Spuj/7frrgJbkxr+f7R7Y8mUU5D/A6A9U2c9DSD49LRNAjj1nodEAY
ouoLtuexjMzFgehX0W5XAEhSGGM/nz42wKK+YOky2ERd0qcXEitCzw7Rf8bFOg8Dwt3mAet0/U3I
Eooc1m+z5lf2dfPFqwRhWhvDkkPNV23Juu7C7B72pRSaD7465lr9s9O779hrHwSnyKnrHmvqnoWX
BSN8mMY1gmYxiZ+JpYMa0GGvq/h4hihxia0bzVyRrXPrFb7EP+4Lmy2O1IcBp+o/Ak28c4+zq1/o
fq9LRpo44lEl5eOH+S8sqlPLbzP6DLI89sF/eyhbFD8u6edjzbDeaYx6SccKGyTCYCw3wd4OD3Hy
++Z/Lql9/rFcH94pD92yfU+j1TE+sXOhP1YfSYlVP2c7701MHs4Q0JRoZXOMogl7fyN77vH/wSKG
VJyIejMDn/VYUjMwiXsPh0ZCln7r+YQFX4e+TwkgI6UQgWNwJ8actjafmCVt4Ub/iLoZf0MaruK+
66HEZmRmnTVfc8ooyvTOIab+4zMULOuvHASfuXEDe8rxFDbOyNe+ED+x+SOijfCooY5DFEZ38B/p
O0TH5rPitR29XK6yMlxC5NTCYlneCpEz9NeOxoOuTMapEOxrRh/CFRP10aakE705DnsVxGBOaybj
LHom7vpjvJKODPFj5SyyAy/O0pHcy6ulJvLUiQuPMvkZLU/vDb/us32ARlEVnX+f4305cWx6+fd/
WDrC3S/JEB0N4xlQL4GYl0WnKMCpnHJ8ofxVe76ebttxynmr5c7QCLVUgVcEwpQCFDHB0rOpEGQq
v6DE5XEufkyeW/bFR8wqt3yw1nUtjIAAY7VB5u4YfpnNSbndr0XZwsrWYv1es57hdWj5DRdZoGwO
UoLV/hsPQQIW3iaK4Ue0xraOEg9+JGpwp0sU1Kn28s0DZPjWZAlKBCkIP2YZ9Vhs0hKr/XsgbPLy
w5m/cAjIBkOYxqNISCx41lNzV9YGkmeJUkJJIQKoRKpmbZe6m2IdsnanP0fnUqvuXBhLnVE8WwiX
fLnlybP2oT7bn7vFlepFsI/xDkURfVQvo/BKVAn10Ve7jOWVjdF1UDwCJxttVBCdewdXxjuZ3u8d
l6GICFdNTXn/S3hTfC1wnvwoUAxA/B4aAGtGLKtkK0gKFPrUAibeYeeYkTLVWnZGoCIwvea9JrM9
ssUJEd2HdY6bh3zbdvkeJqea1vjn8+yicCiIMzVXl7gJQn7jjNR46zqYnVD5x70OZ9L2cS+4pmQf
Nl0z8isdZ789ppOc2u2g9LbaNx5kbK9xfF7fkz+O3+7gBlikdadqcXR3Hfog7RHjZK6TcIobQmZY
7Fcj9+WVQv/mHkHs63b8nEvoBmd9B4gQNm8v6E5UWe9A+/B+2VVoA6EcMHcSGEYy79yM2fnDNTcf
PAV0LoP5vWdVozzpqm8TdEOyKaOnBQ6dlKdgy1iJSXyz1D/H0UcAzkL5AZL2llhVqKAc+nyFfXNy
P20VK/B0OpFjGeOY0we01jLBmreKPzlFhYM686rGad0CXWg6E8elACh9e4i65l3yeRfUqmsPXjw3
iQos3Zuo1Pa7vk+ob+kXwfpM1yg1ItO1tTYA73OYa0X0RCe/70zT1dK84vAWq7jSZVqnHONhwqe2
EMIPXuf+O11OpkmCQIwlqBgFlYxzepwvUVUJrg5dVZMzwP90GVoyE4td9GEzwqHCt0PjnAboXtXG
SNCAwYHVgRpxd1OW+1Suj+hi06q2eEYr3lQuTFVAyHmX1glaE381felg30DVJaiKAazKl3a9k7AI
Vtqwyi1+OeVNR+Jvwzg0l5N1kFoFibAgLCvHYNeEyroR2VMM97ZK+QIqZRGWPkMihflexp1M5hxf
YTrDTRAd+8SPmOgivSdojnr8w1Ytcffb6iF8ljEKQS4hn75Yxb1v0U5SWaagTDAXkRObgwOhsQ/I
TuamJBZ10VHSqgl8lceY0reftv6NaSj7swzIEjMS6BogUxatJ3R158p8IrwtPSCISfe6BGxiSUeL
d7Ra0ZLWBSGQdq6ks3E1DM/Gt+fWZyaccjjEQ59EFMtHIN9fEBvuWKDW+Qaqu4zpPGUv5P4iBDA8
/JdVP/3cIB2wEAGNp0Ant385uw+QhClhk/esvS1B1b1D9uRB/StDxHbPLpWsw5eb9Lsp9NDOT4vF
dhCc9BCSkHHxdo5GfVFW8Tj2adNbgKwoPQs5uNUAU4bGULYOrvxIWaGtvWs7SvvZKXYO7hSuCMaS
FGN9lrALUSjRry9QCMDuupputzMok3we34u4CpBAdu7djziprvcBt7mruBVsAJIemYH0dNckPFng
4ymFAJ9iJMgqLmEzoVtLbyLDs5An6qye+MI6XVdx9AkqxePzVBooWhVhds0+NTCyxqw8zIogHzvo
lSjOFvHQb7MLeVlvKTG0NNsx1uqZjJK4IfMJkgwIw/HwpqCQQzhdDtb1b3wKh8GidgeVqcuA4Nk+
x5Yj12MCP1yLC0ryl8Vym/YjFWiK9ycYRxZfZBqeYFaEKwpsATh3sZU1rulEQKH+d46zNTlDySW1
M3rp5sHYW+56OxAGUfbvIb/0dDSxjOqfeEur2cY29cRe4SKzIY2OMTVaJJ3Iv/nQPWlHjUbkUr5M
6y3/e7mcX81wxESHyfjjL/d//000BKcfaAmrrbZC55U+6gG5aJKm0PppjC8IOhV7eJCw7lw97Qyp
YQWWuWmkgY3AljDL5gIvSeaW/JZhlpmIU+WqhCGcEvxWCKi5h2T/1jQglZJVzPPQnsFo0y9lILDY
uORKFxZ4LIzB7vXiNpUu8ga25naLBeQkSYeV9hkvfIy5Vb8aLM37iTXz0qQs5+2xzUoqbkS4PnTz
mEDsFTL3+f4G/AhIE9WfbTz9L2m5qOJLQB5KIXaPt1e+0XtObrsWfAcqEjf9fhHVVragi0fi/bsq
ic9bd6xctG0xXINwZJv4yrEWDKxe6v95Qc47+sHDjRMt23MZIVE94jT2OjBCEE9CZ4KmGO5JOiKn
LUPoWtI7tny2zkLfeoH0GZV8Lq+NZOPNm/wR+uHKiKXt4M4LDwu80Zgv7QUkXtgFqF98WK80/4Ve
Vlg6cGTcUSkKkud5EcGd7EWaD3Qu6UWcBOX88ITWwPiLMYdX7cQTeWQY5rfk5lDsHoQLVtyo5s5N
7DU++P4yZO5C3ZmmfBMgJNwdzutVVCq5jxInpfffeGpOlx1rJKClHa/WsUhHMyDx1Jc0qXGtfz61
+TJpVG0tRs3oo47OGz9kWJ9usR9UncxJohrc/n0aLgIROflFvp6SKu/Pv9lNJ9bz930PXfjz36ge
+RAaf4UZ+jLOoo/5Ie/xQMhQgy9KY6c6azI1T8xkYTq895C1p9WzCLS5xfMW56gU2f8gtAp0L5CL
hTyYQxDju9/0qW46I+HsNDV16EJrhLZjsD+Fw5x+FmRAgUe3AlYk3eF9Wv65F4sUQJfMG5DyJM8n
u6nxtAmRTp16FEpyQDDYymnsTyA7fUmU2BnKsZBvC89hrnkQ7pCNupt3hsL7AQ+iphlQ4YIzwLyh
s+yX4PWDAB6IMbco7dRPUPVlnKy5WMTreMuWTPFySl/frvUK5aBPYvZXOm1yDm5A0vSWrfheYjS8
IAvLG4Bh/D9btdRzYE7bc2I2/yZptqm1V+qmyGBfJofeFC9B13Ig+4Kn9ngZyNby/b0mEeA8/WoW
Qk/9VhFtCL71iQnJVKjYp3naoExNKnmWRv4yRjtctwLuQGeKzm6zbT4BHmjP3RvHc7GwGuGLBy2c
9/xQnWWOL8+fFlkHxwBnEha9fqEdvyHMiws8BGRUob7K7pj/L2lX5AmPHjfdfRINyWb43arjFLaq
/Uc8JCcMaTC/VNwiU11wWQMepkTfPaJdKz59/7YFjXA2dcSs+AJ9hH0xRf9oO/Lut+F5fP4eHS4h
rGQJunXr+F5YlGpOu0iVBSq8OaJfTSWiGriMKQu5kWfDVHzqQtWShaD3HflhLgCVs34scUXnHLpR
75SP5XquiDs+l2focPrK2jRM21hSXVy94jBN+pM6OlBxR1VujOjO73rKBvvZQlFH3LADgnNiSYQZ
iRhtuDjlWmEllzq8zjje8+GesPY7E3WjWiELICBhPNAZmG+e0NTmVcIELQRsduvpWU796mHpqNP0
DX5kAl9D7jvAEtbcIh0OybKmmml35Qi4aoNXqC0kNmDDB+Huu9CzbnSwYczPX38Md35dEaPGb5pX
6eJpE/2Sxn9dseSGbLhv3oEMGlrqwD4dYnogWsXEDcjpfKhrslQ/SHikz3XA3anrsKmN49+ISiJs
wD+X1f1swwlK07r2PlaryPFHBgHWZjyVTUOSjJw/XnbLpIEMfELIgbcrmzPPdMvvc4CMIgHKYYYK
1lPefL6ubMojh615AYZ4Ny7SVKFOZ/a/u2/kyruxTYJ00lZT4NStEUCMT9mhNY9GtZzgEvrndG9B
2wm9X26GkY5EmXABY9zfbElXqqc2Y1Pk69WTpoc83TTTVj9YlGudVgFSjGExBu8RxFvGaWem8HIy
cu46WOoKdfLMwIp31hR62VFZg0zAd4FYRURbQcHvrDyDIKjgBLbXqhZdQaRbmPgMyPJZgY0YVlXj
vSz1x67AdGwrf06qqH2jKU+yaIDvQCezmP8xQvE22+5eAEOhRJ7Lusfxzu8WKC2IkepxY4MVEVoa
oy2Fi/sQ3ILe3TY80Jxp80stSI7cmRcSZlg4zPj3pkQYpMMecfTjEk/u75pG0sBsck1QNvNC+2ew
/uYjBCQIfxJXqSMTxh9wXpfx2WffhUIxaH2Ogt8cUqQxyKeDzKLcE7bBGs+c1bzHZtCCt8DMnB5f
JaPc1FOQXwWjN76zUYRyQk5nUUX9GhQJ98DKzL0FVyVgeGjAEIE3qmWeCudsZA36c2Y03qgOEQuj
AyELBji3jef/KHmajepRGo6LN88z7fmKKRTQRoAqNe8+hcOL/rdb8Cq3SnXYBmFnIccIZAxauHc7
SC050dZfH8M7jCvP+3UvJKuKtayZJffjnvA+vnb6w9DkiZJhUCUtbhc+m7CefLeFET4BE4VAuRhK
+llXdUToiND4Y2wVquQ25n0AxbpKTXvrQoW4hrT7WddzJXNguNIzlc0UmXdoUucK4WIuUtlKMiir
KErPQXZxwMxsrCMSs4JRhv3PqcpffCrfAd8PVcO1kjgrjeEjUElmd6RwKYrV8nHPWGmWGYl6JR66
u9o8hhCio3Mmpv8lGJjDuUxojG7uev1qtvCyfI0KDWxd7hQTNte+SPUBuqUiGqdsb2kLc1c1eSKL
Gxo/XlfkkpKmMOjWdKyyi3wmZSCV/QqsCENMhK4NfFdGYSp90iP9Ufwy0CoyXw74x0bc8uAQDGyz
1zp6mc3wQqTdfZWKGqjcF/qyZBdt0Q1a3FgZELcWFp/+YrJ7i0DFrOZlM9awui9Eb1dVKdQ/qD/z
WkWiOTStJb+KoeoiCgAZjGc3ZZQrqx2GCTG+kveOhAB5yGsWxaYbVhH0+HrwHOZKKPsYQUAV4wW8
b32q0zsftd/ZNHoI5oVquyt5BeqCzQbPNDalYK8ebUvTIxSH/h/nifU9+sBKZi3FdTAnXIQVrsIB
Ir7NFWc1iRmHyFIgPgsyqFnxgKmr5iobcISH2kBKB33N1F/crSdYAZLYWbPX4znU1x+0r5K1Lo4M
1lNc8m2yyQa4OVEuyD9hXot6iRvENI+aP0Dx7L4mcR3AzvrVJfRyKJjmeHx9ozCK0sIVbsvbXhgT
49E9U6PCYVLdhRritlTI2nBLPSRzjOutAuqo8Y1DmqZC7vgDK0SQGHzu2FmTET+JZXWbjMaqQ4dJ
8ZjWVQQabDVzcJ1vaMjwK6/Qyhug/jiXsFPgCarcy9syBjC+9EoFY9pYHsrrER1RagZf+rexeseJ
b8sJAyZFiT7fdRsR42ChHSFrlAiZLy0C9ToIOi2gWNYGrvoFFndVnpm53Dv3X64707t+9tKrqpd+
8gYsgcORNawjGyWvbB00r2M14y3W0ogZ6IRjZmSs3S4nDbKZVAGNdbiJJd59Bqh2OovumP45IVbD
O5baBvS8Gvt7yyvIH66Z+doSOPyS1d4aAVuxAZoi05Tjac9KZLp8RJVjj7l8ozt+Q5CPyJCB038E
ETZVUW145o6wsv4h8ZAZLnbZCJNwefJWnimy4okvfbExUnyMIS5PoBtzUHPt0gRylB/xBXz9ycMi
IwH7ZTcankhQD9LEhna0ML/8d8frSLJRQs+02dl7MdZOB58kFyG2HzWvPuJhTXLshT/iUU/L7yJ5
h0wjEKLDY1wl5eR91Hrm8mHSsGWbzfvuWG5ypqYBzFaNaUEilv3WXgBH0S4KmK9Qfvv1w0HJjL2k
3H1StiE/UcOJ4sEKwa8A+g627P65z07OY+luMtkJdbQlM+iT/n47iW8SWGYn7dgiS84LDRBNXdNU
d1CDoa+5lIE9YgjMe1ONDzNmOcxx/XcIx8MGvtvnss1Uy8pZRx2Bh5ppNGP+lDAWHDA1jurQebZ8
TVH233/gioPF/1zCoei9+6OoBBLwkBVOirPEJq4PtlFP+/MwTgDwEo3KuSwk1VsJ5FhPHtQWZ4Ut
E66zxVTRbAl5Gj3ZlrFxF7T8GsSqAxrjFruhxDnCM3m/tfJzFfuK+RycUgiIMTI/11dFMoGQo5Z5
nwOKKK0pE0KJIN3N9WIs2J68unRt7D0sM9+A9KFTvfWsujZ6D8zPGNxX1Z9ZmWfUwzBDWQf7EnUR
pDt8tqHSr1mKIYC1n5vbVvlCrEVgchteE6b0gh8uPhywqhGZc0zhw+BJygGLOwibty1LLydunwjp
QfzciZzZq8/UJy0ZXiL/6FcsOuraEyxiMh4PDsw0JzPRoThh8T+OYFbrK1PwvHfIvqdpNCG/ieTG
hcSLOWRC7rRazbsPlCa6jM0zNkwKiZQignW+v3fSRnTM+yF7tcnb/lQ8iqhxjcKuh0wpUem0TGRU
EK4Q5sfbYpuBJRG55THUyXCQyrharGzIl5RLif6l3vM4B8Sm3Z6YR9FElYmXZS3kY800hhJc9GiB
tniks5UJXYhpmS7KedeZjhIBViSia3VqHtFaJa3iNwreE404jnwEfGdeU4qnUWrTdT4RawkH8DN6
1pgv8ezJO+W7HhjiSpD4gPtH5A/NqimYaD881xrxFJ0Gps9bezBc/EPiMWgjkfivqJhLLwWvKGJh
G4ByzBAglF+QH97Mf6wlWqN2oxvwXoMPH9XlM1p03JULmpuWcKsNCUj+v/g+bluoaoBKzkagbfOC
IoeWN4q3wpmPZ+dC/Q+NYUKmz5wUTldO+Dd6WkqEUibHVl0dYfCXw2EeSJmBBpLV9WZ3HqpZBby4
y00PPZ7sK4cjZ4cVHps5IiKG2x3vzH54yHVq3iSAYmkWFREd8zcZEp+CpRbNp81/25FePrNGWbLP
+9s17ATmk0uekHDwrZ0PY2pt+WVUN3wWJmooAyfYmFFvdStHe8alS/w2IwxLuIzyM2gNwSns4G12
zb251dDqRcT2wcuOtogA1kwwroaozBr7d5Hexd5vFNo5bCNGcAiTJwWRu92AiHUPXUasLUPJLzjp
zcOIqIeDVVni+ves0YDq7URlN5kgf/SQKohvlblX4dYyJTExUNQKPWDZDNMp3S5xXR6OjQs5jht8
otS6ZTo8ZR1wszujx70lcvGzXZocGo6DelPctF1Ij/FAX+iuvihWgcOz3Mm+YvlsoW2XZIPOSNBs
eBbX3OPs8lUUqf+KKnU5UbPlb7GBtmchWjUfPSTOvJxbf/EcwZ9CPKNCc12XqE01ax8pAUEZxewf
uhvz0hsVWbX6fJYYUZCz9GjcZq1XRXRgHHz1dpbmSjjuKb/IpE8+SJNxIJ/BZ+cq4zk2vn7XlyzO
JcZqkagWRV4OK+ZtjrozSV/1rv6Cuim2B6q6teUSxoXASXpfslce4VL2AGO7QlZflwFnIwLWRiC8
y8au5SUQP9ns13NW61znxsmiI3GbCjLoI66LHrIjIWu9zoDgcVV3+9gVIkJvXG429YlnmhElO7Gq
5Z0vtDll1flR9r9htQNyBAvXzSz/GFSrVSf/1a+IF2Muk8zfjoxtooaIJnQvoSFyzT/1PyElrgBq
a+PLyMQjHm+iKgEPDqv95W+Yc65T66ma4q2HBzl2NMDhzwmVOBh10ujH0HvfvQPkhTAOCpX0HlRt
ZRTV4crqlZfUMU0okGHlHl84pvt5CgyqH/AdHqIoVUecTuwfILhgrkFFNngJmwP1VZge81Cwk7vF
FOHWVHoVYGFCtRLUDErXzWrzJRQipsxNT33UJsCoEgowyU/YiZC/WaZcELvSgn78jQ4nlHv/iEam
RJ98CI7bVKo+ru4KpnCeStvvSfd4KD3D3QCGjb9Ob9Lq3Q1pTs5Tkd4oeygtjudNsDOb0DRoEYht
NVI+NSmHHeDs5yc7IizFtYeZEnuvT7g8QNbGJsmfyFOiNFaFz/YJr1GGdeLQBcK9/GQxRbwUJ88w
oIiuYqE0qqYrZwSfX/hCVMdv6yLUWHmIt6m3zT/ZGIW3G6b9/HXIFddRiPhTzb0aemuOxgcw5WPu
2k54ZA0dQdCbSQsr6eTVCqw13Apka4QhcyhdATM3jzd2gVHRVR2eDptKL+rrmv47f+xxksPEUgfu
RdmUKhBaAeHhTFFW0sqPoKSfeA9zhPbOy4n2guACqTOFUzT84/dzAf3ngAguB6mNdRNaLrWYvZoD
ZVBT5dhtSaRnPRfnwWyJkmyaG0yboUnDSN7S5wn8LzlEI+c4uMCaEFigfP1gZ6GxQg5RipPxWjnj
33+BPUkn/UD0LZGxMvC5TCReGDjvxIBksnefEoGnotDiXx3Ywh0204YT7ZOMXZpa6N0v6aWckO14
CDkRRPbxgBlSc1WenV94NFF1DBKnT9dXqkBiBl13590+3CdXEaQKLzG0ep8zPu1MJiqkvhBmhkCw
yan4RQZJjDO3iFmnLEntZOctFcdjMKRsh+4AhL6XfE3qxerwiZqWlB4DiEL26pGk43F7wZWTZqEQ
Jru8kj84vwIqhFUsTjy5lUnrlSvliNiGIn/uiuR7OPnbj+ZSqJUj+RE6EppCyVfKZHzkUDYx49Gk
hIf2F0vvY+CjTPctF6XgeMIcwafAGUs+EM1izFAFslhuWvtakjVjXWt4/RSJLhRh0fn9qCGlnICJ
Nb1ktBXUupsWY8rmTt1KEMaHTAxo7R7BepKpJZBY4DbAj2lOtqUwKmeRJFRsDW01AcUGD2qle/Qv
jrgcFHOs74DbCKAALTueruYJd8Gmsqq9KMPaaZewGHrF2Ur82B19EO+oi3ElNDUlhvR0YbyUFj5S
KY2n7LH8PIEocs4hDAHF3Qq2szF5cbZWOghfOcdUcJILyHhWY2zRzudsuQBsbKL24hjv3szn+Zxx
cqo1qG0jfeoviPZIpBNMYIP6Il+TbcU/NzGV9qzPnh6ZeEaLcoqkjARBWpfkum+i8rahx26By/Cp
SYZC8/3lLDsN8PZ4Nmcpt1VQ/BeJm6uY2uVeIa3Lh4Eih/y3tteET1ipZN5dHTP4Mou14OxNmXgT
PqVmPUjbzl2ZlffLQ5VXCm5xbmIS/PxM0KIxBiq94JiO0oOiQdbEMbmYg0LLYZ+7hg7UVHwKPk3P
+/po9hL1vTu+3C+vuMFyeXGnOKLpKQ7XmNxq2M3Af3a6Mj9xoXKYr3OIEScv9TDmZLIfdj664yOa
fOT9TRhO6JW3xptBWfTLxSZdN5UnD6oKWpJXJG0z0nQt4ejcAwVRDB9fl3QcRo1LHEbOFPMUgsK3
7GRjnhoDywlo4s4lmuxbUm9kvqYiYVNgRMajiumStL48Sgv9ylKrjlV1LcEu/h0Qq+hFLvQ6fOZr
srEzyAZd7pbcWSgyCYr3HQ///rJEv/efSrZO5+ewR2XC6xh6hnDPsgWe+74YgZjCAAEZN7ei0bLJ
kRju0RBLh6PN2XCtTcSqitHtDGBE45eDztgSvPFos2rFFuVcQniU5ibju8LTRWxZL6292rmifckj
AfO6wf4R1+/P6H0t4lnHBURWoSaHjR4UQZgSpKwqwsfMX5hR8fcs3mpmMIMD8GTv+OTS6Nvw5Fwi
0+T6jmxhByDTxhc3BzH34rTbF+ruxbqP1qZrsVnV+PphDDtBYYg15SgG40V+Hgdk2smNHxmP7SiQ
aGLybk84KAqnWsi8G9SpZMzHqU46mLo++L5xHXYn02+1slLSjc5CbTsG/0OFseWKFPpAI9S9jIz6
KIIsUhRfpY4QtGfxGAH9aHIABvttVRC805q3OI/l+VwDmMhsytvfUY93HPR3/ScDiJonCSjpaCz0
U1oZB+NIxVVLcsguSbnp8NBJEYCAy87EcO2OxL5VLim01I8Mt/2xaTqGVTsDnDypNiTHSzJbB/qY
pa0nAhFpbp708H9RzqqnScbUYhx9ykPW1uFxVjJnnnebR2prPKjHgTcfzJils/QBTNZodHg8/u09
5z1U4TgivAeXmQMMuVJ4KOOYGVv7IqaYn8udlXnf0Xv6kDXMUlM9BmXNRGuHdjL/RyrPBNLAwV4w
frXH8zGAna+Noa0OxNMPvU+o7CqRdXZodBumo/LaNVWkiPzNDo9nKJasbzzW0DPFx8hcr+bEpeB6
LFd6MG7VKKEKw64OIWHtn3VeGXeBOtc1e9Ucap24Enn1HRfCjyLqCKSaoVcbhr+eGb/oV2ZHTLn9
X7l6y+HALrVLVAZa/MQVy8/ULcY/mpIxUyvCoLt3rR6Lj0ZIoDCs9O6za3r+EGcDUuCe1zqYMOcI
NELZFywmqYPq9CO5TiAlm1BM2lExYIEdaaAnHQGQ4VlZvTFcqzvjYqX9Ty5o+LyMJr0qMc1pZaL2
qkaou4braem/OiZepdKySlerUxO6Q2MMEXilMDMlOiYxVfavvXR70Z1pargQ1yq6icoluyJtkYqp
skeowZzv0zomKUMWjImmwx8OFekgGbQetY3WE+oFeBHJQh+/9IUm5P8lodnMlnxAFiLCbXfrAJlj
90DVHyZoBbD1Zq59PJfMAPYQsS9PxWls/3iv38IO0K6HnNcQbMIB6eQ/Yf8bIcO0DJr0Z4ppPJRb
91O8e8WY0xkCYHfWdE7gFNMvHE2UH0syWtjY5xwMlbNyyjZo+QJa+gXC0jlryej5t0gLe8tDefZl
f+VMlidcdAWYW6m/aZs1DDsNO4j6tEdsm7P4ua5MPtd8wWFXYMsUfe0Q4t+/G/1ZfpmtZ9NZW73f
CWO4MhVIbUCybVdWBGYt936DLfo4CHUVoov6kxdam/dwGL2NI+A6s/rfhSAwPxJMqvzSjvZPRiHX
YdTiWGG5geFdVTAxzq0cJj3t5L80oGr5eg5W+mNIKA/QWOCrNMVYWkaFtMLTXTUfwudDGee8cOKu
APjv0qg31+rNtNT7x4zHXjdbT/mWpxLq1amFRbfaZhOmtbjJ3fpXaEjOEPw6X77r8jh3pwPuvqk7
Fp47HDLGnvJuG8V5NWaFZN86pNBuXUo2VorsTpNnGH0QyWSD2SBxCepLF8k0CXmv47o8bmtbk42N
nSEhtUnuk4hDX19w80+6RmjS8o2B2Bruep3DKIheeWeXtJ6gX5sXGHJYU20HTTJq1w7mOIJb5gXo
k4AlTfY2iRvmjRdXdh2eD7Oe5MFFes1DbqG+LCSzI7xuGQB2KcUQ6ay1IVzmcfrDxKU9KBJRAfX2
71Qtedk9fvLYZk4aIxqhNHimhlJ3YjyUt0OCWwyuY/bYNzxi4F4fO+r6+QM4/weCaze+N9VYPEG6
hg3M/hpfCIetfbScUMpE3HZ7JGiTHNeOmAdT3lwxzICBDxq2fDPm135KU1SBihJRd0yDVTaxDG0U
wIl2fhB+9MbHjfMUh62SY1i3fZ4nM7ERC2rkZm38EOq4vF1vKHBT+JJ138//7wu9cuqhtLMhH+LQ
ApSbYb1InoRdVed/ukSW1lTwgxIUsOo/h+m0l60i+dazaRxpwg0oFxi0PQs7AwHDNek1TB9wPoo4
X/2SOcFoSb4/uriH8SkQzk0NqiPfbprBmVQL+BsX5LL56S+TezF+1yVaHyxtTFLn9UmoRwdYBUJR
Xsy7k0W9g7tFkGvG/2InO+J51kg4yYNr2w3WgE4mghVgm5wL6tD1bb4WkLMOOjFxa3Vufp5qNmTN
SyRIusB7bIMar219C0Hiuqyw3Aasg8OOKDIkFvITlw57vA9rOTLv8+a7CRxVeXMX9zWN6EVrFdJK
efv+no8jk2u5SBAO17vkFk6yLl5s/LzJB5Z7uKAYuEn1JP+7OESWPldFSI86vfKUPuT4wzxJ9GRX
ciq/1HfQ9Pa3FUrkVPcRTwdZ9AmHLbswyOask4p2Uy0P36uHdzHnSMEqBcXp0dOQOJft3DbHQxvz
anej+5vBWsIw2blqrjP67FREWAKyeWjzRTT+rjWlQoZgFtcI6B1vAmbQqk1Up4IO7WobupB/6X+U
8JMGnB1GcIXPxfHMfGbPvNqn1WSlOLDrfHcaIdp3eTzSnoz5ZCC08vvPuwarvvZfbqeyRflQG43s
EP0KzwKNp/JEg2wXyw90pyXOCWSZOnei7aD3W1So4l++zZb1b63kpICPAb2dEDRdirZ6z+g4tGom
U4JCetPThpQT3uvcKpWmDyOycJ+Y7gXBUV0B0IoyGExCvipU63LhNkmXRfBOltJ7TW3bD66BVE3y
Ize0ybbQPqQW1hSqVccJVZA3tkHJ9ZmtsXEr+J1CFfC81sZ2ypXFiWypMTzqAtzLyQV38GFWZmqt
giTIIECCJlVTJy8IaRvBnSy6q3zAEMbCH1cbwcaOicGozRx0oQ1zGNbWUyebWRU+AF0hsPuvnqSI
SUtTkwx+G/WkfMHnjFGJfxpqdqR6bLfvuNha0fefFd2WAHVEFMWMHApc3w8wazNCBwXney6yDDKj
H4564W/LUw3iWEuBYW+QWYygG00pUax8UIJZNqWK4msE7T6vyY1jhJ0h8jJURCtJTIjdTPqZ8iHN
a6xgMwxJjJ8G8a5zUDuUbitFsp2YJE6wksIzAd5un4ZmeNmZRZ1eLzaY4WngnXgYwY3nBQ/q8kKs
FYv2SVY6VvXIqQ8JeYPtxb6F81MXS9BZjMf+T4ILnLLz/x0bEZf9deA7LwqtsyOgWSRlEZTOG6+K
tFMEXPSPPC9vsJB9Y6eboi8fsR8HmQAbwUGDYCjMj6sGLnqxCPJ/zNYK5SOJV29pMCzQg1IH5WA0
sXST5QKvDsIne3EL3t/oFVqcIvIzq5YIIfHGR7x/+ADsLvRQJ5BIrmQPOOV5VlpZSSIHmviuZIVt
aJR7mgpaBVSdXjyW/ZnbFc/9DboioAWpuacHb8fedhh2KjuUHbNGMxwCoFjvStmqARhAxys3u5yK
R5qduc7EKX5H+HxiIr7ZkblPvSFMj/+IVQAkO2gZZqbanDfFjyjCkHqZ5s38FpGQ1Pbar1THMTYG
KSOehDC8VV2IiXGqRPgxGDUOSgcpCjnDWjrfiitu2/sgmhkyB/43QJEYVwNgmcBrNlPj+kvW/UMs
jjWiGvZhpdBHBpgsKixgy81zWtxLtqbmZfNeDDCEzYNF9IgYrTQ2mhzhi5ICz5qvx1c4md87uunk
c6wHpiNCbKJBuKhnl4dXyeEB3jmFiXCa5nYLXfRr+qrB3e4vxTZGNqlFA0TPIaN2aZbDkB7zHfOR
x3NC8PdxRCUTL3p55pIZTWtAggF9WBq6nHctgd1qYSEcAMmh+cRk5RoDf54l4nVREnAf0zq2F9vr
Z9HZvhmzA8BecLRzzI+inv2CjXnMCFHQOTXeNRKMD1UwC6S2E7rA2KctZy/bI9EGamMxx1FOFc27
yQFanEFOxVPUxy8qrOEwFgMt+ILgka4AP+fz9/GiWw4yoB6RK3RCzGlXxfpElbDpasC6ujlBJ0G3
Ml0TtTygrrLPwebo1N8XhuIehgMerCLsS3uHCUDNrbYyvAVNavpZABPVHQFMTo1awV9fDBNA7ciB
QFKZCnA/4h2OxNMbbrDXBhOPFAP6EBrAf99RYFLMOLhOzJCCAmWJCG74R4gpPb6klUAmlawbadv/
16Q/Pi+d2dmatvsmZajQHNVND6o7fOtF+HZrSzQ+V7LzNQ2lvbwG6Jql4BgFNSe4G2rmM52DVq8A
LA3UT0/SHpZrPuAluSl2gtGiviO21rhNP2rTwyU6cbZpy6heduhwqyR23NBlRF123+2cSxzXYPU1
y0aaWRBUWqs/uj7Gp1XGBvpOeZKYZrZoVb3LCdeFWypkTpASspjtA545in+i8RQZV1cFPNnT72d0
sSYjarBxu0IIBIASKnTSgih6gyzboIfoXFplJEjMoJ6xaTS1dI/RTdgH4s44O9l1JuMnQSgMe4HM
DDBMH52rU0Mxm74BMhlQlStHGP850xtQaVURX2bAfIobDGzR/CDuLsHim0i2g/zwIc+NJv8hYUdF
hPjeMmEM8cNjgIbZui5ENQaAeVAvlIWalQG/pDW3Krn63UBtqYzCavd9ukKl3GDU7H+bxqt8Jucu
7KSzLpnuBqMfVrf+wwdsYJ3P48+W59Sy1lfxVzgips9Z180agbxFrdx3UbQaT4Y9T8051nC1qYKf
PdclkX1PDu6cIij83xCQ0Z5tWRmQAAIuTOcbI1FtzsBB2+oVU/zGf8sJB2rv+4+eh2ZqVCUY6IAr
zqylJSHigEf+FI1WkjPeyPmF6Ino2VrNJE2Rzz1a+pjMdleCXJGHfge6s7YxCkhROTaHM6TgOz66
5D0/2qSH7KFdUN8XM89DuUyBRs7TvFa2dInBBQR5VdpynqH3E2c/t4bRVdnXfFkCAShLkAg+as2g
6QsRPF855N7DyINK3Eg6iqVnwnUAD5akyVEQrmVtuTUOrXqh8h2qXG6WYbew3OpHBPsqOqD7DdQL
qX/wY96JUGvoep3ovoRkzP/zDK+4WcrUh9VnIJozQFhRjHzWnK+viO/3aZj3iTvwicOwtwxNGa5o
/7lERqtRfhYwkrORoaynap4w2kcZ/FAuCLFapsHNf4GTJXZbfcKjAcLRuaNaaju/BZbfgTdu5lmr
O5aj6uzfDk/CMKOJ7JZ93lHmi/tf08wtOdNFnJpaPkyYC8iKw44+AmYk+UJHcjIvGjmwEklxy710
KU5ZGL9NvZ0SyODF8e6Xa8wbaQmSi+fvj1lHbDOFIGizKjw99OEiPmaOZqKejhUv5BQHuodewCN+
LC7IQId76+Zu77c5bB2nPZXe0BV47350De9Iaf0poEwFqsVL53TZJvtMKL1I8ER+xk8NeEVYJmsp
CrvXjgjGodwMBWki0rLI9PBPNjqe9qTYH/OWLHWYWdenuwEj0yfajSEW8JGvwLvbJ21m1NXaKh/a
Tb7HO0GzWfb0N0Gbkcgz4ZXUPjL7P6MpGg30ACPvyXvYy/u7T1OLkzbVHXSqvJUZXoomTktqGv/w
le4GzlFxTDEu6H/nlgWmQ+eTH0fEJ5PTnL+w3QoUFeD2WaAIEtZxHPOaaonSA00VyBiPZMfAhkjo
BmU4B4QDnY15RCf6Bv8jxM5MptIQsxBDRa+d+/uo5V79JFBgBJQ273OQoPrBeQCMFszI0d93WiGE
+kuk0H/YkCocozmzsE8QFKwdk9bsXC8llG+gkUi7HFApVQimJkJBuPpliypJHbteixjmHSUN0pkh
RE5xiP8qHGYzifOdz/CBivh+J55lDzCsZPJXfuQMgucytr0Ytx+3UnptbcQCMtG+JQHrwQ5f77IL
KG5Wcz1Gh0yUhdZlwpqDpVqYbGeKx9d742oldCXDTYQhKtQVsP1T6upmoSxWSyHm5QehsdAEqpP3
vffLaFSH2OAAP1Xe6QZjDexRd2qWoSRW7e4u2qmy5wNNKD38vhBVncWa7wxRN04rDun9UiKCPSLU
hrBtwspQi2/C4YtGYSG7gc4uJFLwY3HRasbkADmsBVUc3N8LvKC8T62Ot7/xOYxw54dgp8dDn1KL
NxT90to3cr1inf8NSR/lV9cqCBoohRubx5MpxipvVFParSrQlPAiFjiJiXHQ88HW5t0CDgOdQkJP
zDbZOLRvEb8hVCAxi+9EZdFpnM74Bpj31Wup1/pnkwG5ierMW4JxeS3WX3iUH40budX6P4IiZe4Y
thuxtqbEWo1r/fOmYHsF13XodIEW2xLZenO6aamT06MPt9T/ncLP29GxB6xfGAH+xIi2QxUI+2ct
LGspUmFZ9HwJqchNIuqdN2hnZ61YZnV6P/CE+cPzcMbb2ndOUigOo/k4YYFwttDiVM8RvKopPsd8
YwfqUcK662mkaykAe6RhAk8uArBDJc9TX4CTdF/eaJFDOzFW6rWAgsYwHwd0MTXTOnmqqQSY9T0W
Aw3PUT/AI3m64RQ1S+Nz9I0xvC4Me5YsbNe74FP+FY+e21Agcoha9gwW3qQzUlne8uDxAKwijc6S
YMsQtLbXG59qwuhTsZOTMN2c19Zzx8/nuBuVC69zpOEXUCbTbPG7VoJqF+zwIAz/GL+acU7vusfI
P1thsy8AXSfyqqWNveIGfZZwzpWB83W7rjXMW9UxbTUFmlsxWo4zJTtiXaCMdaTX0GkDcTdddyFH
dMJus9XNhC/j7y7oup4nALckt2c4Nv8rwmStVt7uRgsWzzcWT4ti5Vh2F8kbW0OQ5EpawhKmFdCy
qZK84K+OnXO7Akdp6Yx55OxTWktiKeHPj3cgv+jxZi4dDtyxPKXKA6a0vTyKvaP+2YkjgVLxVZNr
1HKp1HQ1fx85PPGphA/TrROVTBMKHmSKpfMQiP38jFqtELgM8/8pwaUsYnu5e5e2wb30FU4PoGx3
FLh0LLKbplbiBAVWw0aFZSY+sUc/1n+T423FoYUFFO1DsnSxWdTkEkgnulG9oMiszS7EgCr+sBAt
j1kkbAG1IicbJsaY0Aq37Hkd+c+mtAYa/lDEajUtuoqs/hVW6TrjYZOAgQE92Q5o3x4QFD6FlDLn
Rj1K+FtKNTLpgE8R9QNHjKpE9J4VfBQPmcw8HJD6bqj6vBMllxF6fHknweRdki3qMHjIISopFfDY
VznFVR8Cxt1cMxTF2tSDBm7Er/jxXP2Gr/bhlUmxajpk1U91zM/4zRQkzZOuoE6SN4lyaHUzNM7X
j+D74QVv5XSsfNdQfrqNNXNsr7Kg3AvqFOqaisAC66ULT54QGFWPOOpLHaMJrwdFtBjAwMoAJybt
87dwCk2OUkpaIoUH2VzhhSNhnyVDwFtc+qygHjNZEmsFwfZlfgyF4wERNOmpOhx6xsKQDazkPL0t
VuKaScrCi2LzVa17wCPJbyMN/FnuI7WSrFBFmiyNc6l8CPt25oeYli+Nx0bzhbUIcRRA+lbTcCj2
sPC3rVRbmc6ph5ksrHkpKaX1tz/mihCvyUDLZvgom55+i0dyBohEQIT16/g5SpzvSi726B0CnQf8
SfGy6FCSEhZRoscLg5XS8HcQTP64wtepPg80JQJIp8wXEFP24uNNKiQnUZHcA7yjWkaBFloln0Lz
5irAEE3/tQvdPSdrQB9aUrwO/aD7HgQO0yvKVHN2n4z4OljeI0R4ClfA7XaR8674xS+NWj/TYFdT
XS9sH7jH5I5rGPc7XrlDO+eq0aH+A7ISTv6SgffVpQKiWDOooLIWybN+qMkU+DiW0/sPx9voDOtk
1wlkVyBdjz74sAWtnvtymVLvEk+kwVL1P92uxsMskANa4pT0Tseb1HGSPPWZkT3Ml9hbji5hVyLM
hDMBwrvEShVw/1DijCTSKLM18b7FMJnbsB9qXXUU043IHOD037zBPJGygFEzRUIMiCqSUdGsNR48
2rNMBiuSquw+JabKYJmK/cF+nuTUuK4EWys2dpP284V1s02TjmebgNLi/M60/mDKSP8Pt+Q5JdqI
vQYyeIdu/h4B7h5hbcoic9zo9OZKic/pgTtrSkIfzsjQG2rQM2rd8THVZZL3nzFGP/B6zMyrzrQv
TenbscGx+GgTbT9NvNGMDCDkqeHy7M9jojycGsCkVcrhLX+1pWxFRAOiWYyZkXK5PYyPS1P5doNz
IWt2xh5THEiqRhtJwIdBcdWIQEQqYeBXUinfDPsQBHS4ReS1D47TrVglsr+K09YCBHRELC4odZW2
AHDqnfEreyky7wA3B2rzeHKdxR5gHcEDoURy2EWmSiyHUzM/4856AhmLnTP7yCnEJinhoubS06co
bD0y2bqtKPUTzmvbZNymMYpV7wuUwaB5zVhg8IIqDEbX8DcUjCXf3ZjbrXHIoWNvpSNMv2We8+hm
0LAWWRU/gW43ycomDf+YhKfs0++zVf078puTPzFLTZdAN/o5fj2TA8iUgf0kgUIdFJYAoJYhg9V6
lU3gAlCfB4Lv09KVTCG14QnaBlrrmtKKFAn4PJbGaznviRYgrszOb4jGbrGaI6sMPuj4RWkAFx/a
JfaqnX12tyDqHXZnXqJlsBvhXiW4m7iwjOn0TWLADHcWnvdBFKG9Fmd3UTHq0qswssB0zx3X2G19
9uO4C+j2NdZqkAExLrq4E4MrjhCWhKPmAi8/JfjJsGtmEOMVYfGwXjooxX2rNRnhfMMhUncjaPjS
xGuoIgyNXoUPtuDwOlZ5iikpzwY+Z4V9kAPlWO/DqY6I/snBgJFbuaSyPAw1Wb3PD2fN+7ucA77h
GbO6GdUo9dzyN0x/S0/HhNxXPW8a8iQd0ntAL69vo2t+ddJGGW1p4pZ4g5gqon3kujnD3IuwExY6
JMhKCJcyszfszRA5DyrucpqudRkEX3RlETDEyXrgs+RVlkIJmMJKnizp6nAJdQyefmVla8zeV3/0
zzB/kM6QxyCbRvO4RFOXkFgjiCpA+5Bsfb3X4cxi4KHntinM6K0M1S93rUewssuYvP/SpCmQ1gxx
WjOz82QFGwg3zbHH4ffEWYcrnVzBlmnH7IR1SQHrk4Jiwd/vAgxz+0OGWms8BgOBZPpTLvEgqm1F
k2x31cjWNXpOMDkAJsScXZJ1h7LNG5ozIUE9tRW1F+TPdKdEOtJwJUuPP/CP0L2GC05cEjXgW8fO
NXO51iFMRC1bTJmt825YzYWEQhufAWRy32D++c+HJrZi5OI4ohub4EiNdSkCl9B5VqKDDUzVsCXT
/G6BFhDg6kxwa9WsLsqc5o0hkFsNlUSUWlUXX+cToO7zVQWUDp5Si0G36MYyBC8dphESCub/nof1
HXDm8e2NWQ5I+NoO3DarqKdMbc9iJ3RgI/y4R8cfxMacuGdD9WtoWxfBg4Ysb/u/fNwc5tKF7Q95
mJ+C1R/YWHRyQPp2XbQ5Rg5ApUdr/OzHu2ZQ4fyLcH1MbTWiLljwP9gm0aZVjLwnNcW1vNmqzIFa
oOCcE9EhcH5x3Z7GzUnjoBI2Wn0U2ufJk/2iWuzNQkb4pU2VAqs+DMwQYPNqYrBcRQCCbvae3YKV
MPrhBOla4zFhxezzocj3W1iNBdFiai37iLagQkb3QSLM/0XZ5MU3oZauNWmrhJL/gIfhd2vlyqFK
tLLmcMEPbU31WtpdEHbKf+w/ko9PQmjnIbtMnBU33yBNrHftNjPi77FuLTGwZP2yTBv6Wmz7AR8+
dc7U4MbyXDvGOdkH1fgKElW2/fBgcrlqMtXRQqVORpNIFojE2J3jWSX056IN0j9Cs9ACaCdwnP23
bceUGWVylPtuuCgmyu8nOmFUCzloVnkj9jPkyqBLcaK0qE+GED2QW7HNu9udUsrdiF0HBM73oNFl
0NQasmtbCIWL/OL1aGQJLwh3eCyUaHOTAsSVuMIZz+Kg76kC5YiqXEySWIWvggjUqwqnuYrIWwHd
pGbpn4ktQlwW03gH3zsVo7Y+BlTZ/UOl5lVlOT/8/m+IDgmGz4X3m+iaIHLHO7oINp6JOYolTXKs
EudKb+wPHAUODBbM5lBiJndljF6Om2cPO1+Adz7kYEMQ80xIOhZJ1wsVd3ibIv3AaRCrBDj6Kw0U
BTEZr9ftllXB1oUn7JhBLp2JbRj3A1xlv/sH8rPy/33gub8lhRHPDkJF6ZIznjDNlf5oPZ9d1pSY
ovbR6JOIJlNSDG/dQDsd4+QTC0KxNuYekAfuDzevCkYkcjV6xh84Ieg3lTjHVSUh/C8aMA5LhBdX
GfHBqZCx+RWVUbpvY2ad+yZ/kmgaucqCGOLDfDaVJ2/EybHP5WABdXnDR/Ot2WRu+vbgNK6CcFT2
9wf4d3JJk3kbq4TlABjYK5HYu+GYaVeqGrj9/bvwhrNYS3n0forSgc4TJ/v9gvkEqKkX1o9jLM30
gEdpqpAb7HWEWI3djtUabRBwNHXzU3m6Ku+B5cgKBNzCH36ZsJ6FHUC7PeasPq6a5kvMCO2LB6OX
SmVvRIz8B39vNthpcW43PUi48oFpDLsL/4dX7yadIQjQxC303wI4Yk2d6ZM+AVsJvE/VmpBlCyAz
wzPzMDS146fzPSTEJ7mu6zw6dOuYvIjYSITuQAhr0Adnw349QQCLxLIZeG8VdSXkg1R8JolcUfdI
o+4552OQqaZDXMHhtkfSTxi6iF2uBnavdQwrYxQix0GMbxGoNVq4f/5kzK0RwBourujYFO8q97QT
tk1VGCNJxf+/uvHa50mdNlHJjOgmQfNwwC1npUmKn37zJDGIj3tBpB3nmv3d3szNasPsB2ORX+1d
Gq4A5orp4iMaNCqXvYSiQM1WHbwVn+BfvZb8VP3iTBwScY3S3j4ojMw7sFdXPBP4Q+Vs5laQkk9s
NIM/uAanLKBtba4wqkQef+v31SI4BJOmLW/JGk25WhO/w/MqAAM0I1GOr7TE8QKTf5KjdROkQfcM
LDoRjnFCYcZYmVLrna3/0VG1rDipgSRvL2JchLnv+3BnO7sakKKl0bhIlz3Ebx5Y/WB5wOrzE+mP
omFf6dKnp5A12TsJ2AV52lnNKWtsjWdjhCyJpxoJKDFftFeOXEDTr3CG+5nK6MC8r8jyK9bA/yof
Bn3jT/CggA9VexXYEFO2AEEEwBVaniwMQOn4teRYlOmrqJpJHOEgzcnlUTnjZNMSf5ALj4emVeES
wIDu0lVaCh8KccZor6a/nJSYeMSV/ewl0p08Pek9R28iYEcs6e8R9vJoiERLe8VZA84X72QbzTj0
9CvwTV++nR8Dsb+7xB8nx5X/PSdbBl0PS60YGKpJHlF7qeo2RRp0e61FbF/T+Rr9liKxBBRtT2vH
FTL3Ke3I7ip368M7a9n7VZ6cNgAm7ilkWMRk66pwNG0OCfWFnYhxj4DYTj3PEOwMX7uYci1MR3AT
XAHUZoe3BPLGVRKz22glXKM/HT5EAmSXaS7UpCnCFqB2km2nQFgJyjRub+ieCqEBwJZbt/ksqEak
yoplylp1m/IYz03d1RODE+kjKtjSUwmCNGq6b/8XsOEiRzH5E0xeZPAOM1IlExtMjfewL2YaCk9G
j6Jnr3rA6m3Bn8UVVO9pver9Oh7gd8T4Z+FNaWimCv8lnL1LTNj9eUOD4PFaqzzRiQBoBWsq9B6Z
ZD76cusc8za8Wqp+qwTfwihcHgRV9UjWn0p4e2okqY5Pmj+qPN2mjq+477RE1JyLBUbHO8ElBqLc
kejmd/RSb7hAi/Nuls9mEcvdQ7H8yDgziUNB2fukPOAksFWSXPoBWuNegV9Jw7ShdDqwqk+Wi5P9
qrRHjJh6/a9h3U+8AZ3eLozNe7veYqIiQGpRdRs3WX2hrZGuoPvzKCwwyOLa7XgCXZZt78oaFnq7
5bS+qKS/oxr7sUsRawfpcse+fICpfJUEA1gnTgPFZd2uQrvvgqx9wghbN75zIoNX8RvvA3C1oSul
hAFvb/J544d+HqSrgR6lmEzeRAxvOxR059ztaQDOc4xk8qpWmRfyGQS2DVJTmh6OPsuU2/vwr8al
shskQHQ2GwDMhnn2sB5N1ESMlXkhwzwHS50+ojArENhm4ZnNHit8vyR3vdP2XD2vfXLuABZJ2zus
h4u1+I9Phj0Z/BLK3PYRVsk3wG2j6VlOwJfcIJMjLuKG6TvKYUapUk6riS2Ka8TxeE+YibrJuYb+
fOkNNEC/8uPlozNEHLFf5jWiHpXcLVv+/eRY+SkkXqfekbyEWbJMBpaq+UJnG4nHBa3bL82rIVr+
n+Nt+N7JaockCjwFTfwuoCRg1YpBgNzW//S6TmSQC0dC3l4NDbg6+pgLKE+Enda8zunvnpBkM94P
En+ZqQE7n1d+7GTTYaJg1sZ1MnNmm3PGAFI8KBqyzYotpSKiGaOSzopdp2FvLSSuI2dMVhoeh3w+
+zd1TQPuFnYD0dERTKiw093zGzY0NhQ08FPP7lBPekTGe1dDPTQFecAqJZmkk6VJgF4dhOo9n11g
fTg9NsGQmD9tBppYpWCEl1NxtfIptg8OYwRfjfHkFkHRlFHd0eo7cUxh+hu4YAYDwvxBfPVPvqh8
2YloK/IQLzjuUwK5VOczwB6TzWXM63lqVsHkQkKu3PWXHfO6gkaHEl/F+xNP/nBTE2Tt0Q+kwAVG
SytbYJsW0/uEpCVQ3VjORW8VDx+B/CrOBVF8500Fmp1VyLBbVEfJ+e8P0vE8YnE2LRPgZpDow+pA
6SQUrBScOuqp6qZgcBBCZb1MxYLa4FbE1ZBZ1l+x7p+KR2O+sKmbLmRi/DvqYsRiDdzxVarM6jaw
Zt/eDlUpfF+f6uqjaNB4U+26QO66YIoto4Y3/d3/CzEKaw+PzJYDQt3Dp98bMqM7XsPceulh0dk3
kid8yBuwHJ5nT3MLrkCgkLr8vyvB5DiEvw8LPzqzo5TrBqM7ik8U1owrjFR+46PTpOZmcaVIBRGH
v/eRBHYaa4oJPm0J0nBFWFYeYHxNz5yeWVnj3sR63hJwW+0YdspNDtkT6heQFYmQndKa3HC3m85O
NSerhZd4NYiRuJEkxcJtCEscw41bVMtBKHu4xz1VpYaTCKTuB2yLK6HNFpDgtxrUyA6VWzbfJyB3
uNO4DqYrVe7SF4y6YIGwOJapRQQ0EzwhQ50ba0k2Bh4jKWilP+RZpX4Qonusr4UU4xDav8nsDv05
X3fruCBdpv+pdq7FWpksMAnmSma28pm97oYW7vb78/UNwv2+hjoEda8ICusV2MiqKsXzTTxbQ1GK
mGrG6IyhZosxrxvY2D5WSIb4L9i2vWUcNuuWDzR3Csw1exRbYNKiEF9UWYXprLjauyOfWmWbozya
Z/dAgBiAxqWpgUB8U/7Z+FjBZkSAIutk03FYMk3FoRT5Oo7UhggHtsyb4UsofF4lpOj+cMXY6IA7
5U3+NS9ogYMjcbfj5Z7Jkl6lRcx8b6qWr7dQ8EGpAaXyO9GJf0wT3ObK92oGpi6GcEJKjKe0w+fc
YbjaRrmEzCkOzHCWuLHmV4dw8liAZhZNQQ/kXGDgameLwfyUSkEDeEyPpPYJHbotvyckYGsTL+sK
ggSz/e2KQx2HnlP3wMQenNfSGI2TzCZTSTE33R1nV3oQ6v60dKPoqgCsuIgTSargwwGdo32nND4a
n/1e5OS9MtzUkymsGzZHoVyiQP1+Ot3uaOsFgoGA4bqCtAZW/Hl441IipSBpTPLf2/1ioTIEpDZn
uB3dzBE5tsre5qs2OACUseP+WhGZ/4UKCloUprkzZc2/EQjbUivduwQzH6iEe2TW66VakM4+pu2S
63HbvFXwqgE6/sPGwPLwktJbO8CnVySaPIf0198s6DgSPtVjC90UByPDkE6Pi6QQtwWfcHRl9KZm
/ZAXOYBAH8/ZqAcYeDGn4mNWtYGRecYHZHwRTiqblIRONIaEiXfABZ33D1XEutYc3Xov2tcbGmWR
8bs9D6ZlPSoHx5bfPC5HIjv9EoXKDN9BpKLjfI0QJ+Pzqo3KQBYQth7lYnxfj+ZQtp3YUQIutarZ
Ttl/2YFiwI2xbFDBVIIo1dXCCZLmqaf0HzKfXopeaskfJl6QDy9/bGzcDnoctOjwQ8gEc16GObVz
Dmjh0iukBaVTC0LomhYMERNZ3ivz4gPFUMLrc5RsOnE1mBfVDKW+lDdvETv6jbXdBEeCR3BrMOhk
wUMeaJtthWzta5mynPsZW/uzpz8gWr/BNDp2dCXbK8sPRGrvysrpS+gYf+W5aP8nOAuAN7fQtZBs
fC+2uJNwsg4101/sBP/RbpfGzSOFzyT1RaHvfgHuHsAd85XUKjfxFpab0wFamJBHCdczXV2Ia47U
d1ysV7H36RLnxCBsaCxjkfb8CfRZJB4OtppCNHo6hhuRJVoV1DiynTnJ0tv3+NfcKdKKE5lCe0Sf
0WtFt8SqiNoJrTDYHIq2iOlOSvNdBb5A5PguhI+/jzJD9/mFfj/uliUMkeTrSH3mZ4HX3GLSgclx
j+SPmHFVzeFjm6+A3M6Xi/EHy9GRNRG4rfQe6OFuLGc6ry/wkec1eFBRjCKY8bXualIAFcJ2vdcr
A4j1bAxHhB53jSe4/DK3eEaCP2g2phHdim0gWLYpVatMMTPiLZa2k59ev5Q4Rv0cArzvlyH9skX6
04mzNAP3OoyRBN+kJrAmmMuBI5dgl0Rr0LP/EQqkQpJSdJfR2p6VRfFvpaF7hcrX5tt5H3S2xD0Q
L5/DSuFhiukc6nWQIjcEazh31aX1QpkEBn4K8axd9c/CWKKR1mChySqlqY4NbxLbk53FzrgEaebZ
XV1uAu+Ii+Qgzis22U9MiwoAklxYFIZZNDXgM8eouvCAPkDJDRfjTxUAC9dq3QWd8Yd3bz4IPoFm
AUP0qdmtqLpGPk4lr8kmqNM3Bcd2eAjuW3YbLuy70MbMDVF6uG2sjEz+8v1CNR4ObveZYP+n0QXE
ycB/ay4HLW4XKcNAbkJj8f0KA4hGLVjP8FXKB6Z/QALei27xOPgOWossZpOH+MMlKtxuLYbjrv+s
EIv14D3ItSZ2CaoGorAIe1UarR59r5fdK+2VM1MZVMxLMhaWATS+qxU/Tme86K7dK1xDfrJqUggX
egh+HkZQbBa/Fuxt9DWDc7OB2tv7U9gKonamuj+AvIkROxKHZrSQc5aENUFtWFdbku4hOflzAFcr
Q4RKgUcE365GAa7PA03NYjZNm2IOIXdmU2d3DkCXe0l/cJ4WCm0zYnbUzUnQJhjTm66QeCfw2iuA
S5QiDnrMCJUUFTSmYLZoNWrXVfGKCcA9QRzY4CiIDWMPeiOJw0Ja4PXAe4GwlSgBgDx/D8YtQ8lO
OYgl38HixYSIKF4Q/Ne3+MBd1GPcfRkfUJIpNlIpzf1MRWv2OzW6hPl6k9uT/9oFH+PIZHZ1IpAR
JQwk4rIUMmu2au3LdOcP4VwpuGJjJAvog21HXwHyymZX5FC2lwDzCaRl2B78S1DTm6V0kN/I6qjh
MNgchYliszyUWRWsdkE2NZMLyHkUM9mN0ZyMBqLl/zuZ/TtH1dmOAwk/l8excaR+mqYYDqQGTy8m
//fjiqjBPjkIOjRjTrKakIuzL4YXNHKw5OP0on8HD0Cxg9dgjBE5naIoba2CxjFAN2bZBEtRuSHQ
7EFLf1FVZLWAJAHPxncveFVG5402B0ayzNPgtj1OMGtaU3ZAS4zaF2nLLv6oempaCwNw5ejSPRQF
7cV/SClBoc669+Y/RNVdxlkmDB6eoaWayBOYspD9yawz74tN8bq7gkGgEZTarAN1qFU3h/6A2yLA
ab/6nUyOUJg2ihfb8BTmhFNmRttv1yFkmFCeuvVGX3b5oshsgpEq8dxr21y9GwNyljsx6rqU3Gq4
6/7uLf835HYbfkc0oavDnZN+SnAyMMkKFiTbjqOcJWF5p0PPtfRCt/zY+DgvMTDlYlamw5k3h+aJ
vpJV6ddA/BvW/ZZfKEAwggY/ukQe1tdw1jzImzyWFNFPTYjKZvgaVrnHzES7XQpofq0rFrPbOwyo
Q0PnJGw2yCXOxtRG816nB0Y4Lz06JzDSOh6npp+fxP/x0HmcTbT2zY0AAZJewAD0lITyCC1pDtdn
/5dV0NqXKEijpxsbPaSI/3tjpoQubE1uU1B0gQKPqnKPqohtFFahKCucH+iLaUp/H6G7anxw2oSl
vOxGIbFLUqChC7cJ2E18x0ydLMvtIdM30gqfjvRhxrBWefWVUpjyFmvNPOJ1zYMKEQ4NFgHcrkXQ
tgNhLTdQWvuyknGuaaggMzWwielRUPiKyVBsl5kY0yUowB+1eglwYEjj5wrz8toj7TsSIbGFhAp4
QQuR2ZftiGHQ5qmx1AiWzdC92oJArv22CjNcRkOSl5xPW3WoawbYz9YY9p9QyEFhDSiF01JnPNb9
aU5u465n2uwZ6TKgGjPjc1s23TNe6Kiy0JsSgqYVH9M0iC8tE2+guZOvoiva2uDOLeKyIBi5lsT5
pyT+6KlqyPJYcv6S6oK9cG1QhB//7cP3hlemp8lDdhtAgvbZq9IpqP4k/TVvPoD3VtwGffxo3KCO
6FwKBOumE/4zGsZAdWY0GtpuB8UbH+d8Mc8GEThnUEdinM/+CfiZfL8yikE1XUwon2W33yEZzugB
kaKkeahS1o/1lOu9nzi4wdx+Mu8KAbfKkL/jJ9yep97gm/kKwuM8moknsZA1yFxxhoSGn6PCQVcT
1Fr6Ju2Kagi4U1XY
`pragma protect end_protected
