// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
klJZ9Wapo1Lbe3eXmzOXN2hziBQ2zjlj/hd622lRp7V6J8Z6YZyndNS1UGLgKM66LH90/T5V8/v5
ce1kkd7VP3i68jZS8u2/3uxNEY3RDKtjJz0M+bCx9uzc+FOmSB5/rVwkhp2p3F0CGLjnFlow4BRW
5C7L1MO5oYERHLIH6R2K1H5PgOUCrRK38tEHzgppZ62HYHtFjU6W/LGtY2r7ukygsYI3lzz33mWN
ZyyYmUL5gCfx3gWamWn+d10T23nB3kSq9s189g/Y3jwrWrHMUmivLlMAdsroklin+t0BIes88QxD
P1/nPKhhiCozrbekKF+YEm34NPxmayM35IlShg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
2yeMNw8GMXT+m2P8pcZElamfGV0XVm4EQLY292nC8RR0GNjymZTEYjokFpeNsM740wID3ddUNeJh
B4+4n7+zFWmMSYR95qlhsTUxk0Dz+kW82VejKDLng+8zfU3j7uCrrOwh3ZQcigcxj/n1RncPQKYi
hvcdi5fuT7XatLU63svmyk9pPZXRZW+s71UFFWo2JZXp5E3dBjy3i+MdJ7IqwnYGSUTs11o3UHbG
Krg7f9c+n45pYU4tupRcWfexuax0J12fPGvhfp/YxoekglBhPoduz2lAzvD6S+6TKuAXe1k1b9TH
KfbFmHs8aNfiKhCqWIvacR7+ci6mqAf5TJVgfOubDejNS7puPQZALLmpIjU6N/50PZ6V+argSeci
NpIs9yRtRQvfYUWfvQ3qq4V6Y/SChk79eZONW2G/zsm4RIK6//qCfC52I2kPska30MdUE9GpZgWD
RE2ukUAoXMXSD6g64Sy1KkYOp1I7L4f87t3uEElvMpFyTtweKKpynlopspmyrROmN7UTxFdCVjzZ
1BEdHrkqnjOnwM0lQRePPCZmGiy4bhbh43yWNizOsOAf7vIgpomSbF/2uX9rcoP89Fh4GQ4W4Zuu
YxPrbZwuz35osktop0IV5VpTbS3iNMexMj0rRsLdtthGFMI20utDSijSrApPl3N8J3cNP2u5g7cD
nFBLTJtNYlRmD2sLbg/E/AoDfS1gzPXJHCQNMqKQW0qe6AohXoeLwt9KMo7BIZTiRhjRl02vMccw
Vv0vpLq0dpMmZEboP3FGeJcP9qfrKn8nJVcUjUDb7gxtEmAIkvCqAXf0ueggY887bpRL/VeTVn83
joIQFp6pFzzib8pX/a7hNx3wB0fz0+MK0oCzCY87hV8DMbtF7h0TISjL0H7+AU3MAbgryM4geXdW
8blrGNXxcX648ErDhhoEY+mr8/ro4rGetvO3pWq4O7mt2IxlebJlq5okdOQJFwde1tC0yWOpmKkB
vVO0SWfzi+NXRJAK55VQTTnP+ZllzcaEKZIKs8j9JPtQLRayUfPAd1dkoffsq3Q4bz3PKlAbyxEE
gsUxwPFE14+qdc3r6pM8LvhIFEG2Ht4vApeuGTbIML5/TMDpMbGL58nxsXvJ4WbNrSScfWJ4m818
OwOc4vNorID8vfKryIVz/kyY088IMlW+Xz5D/AUwqx1+1t3nEyrOi6fGKAfzOnr4j3gypc+gsEn/
yd6pLjp1tPvVajId40zkFJUkCcfrLHnQbgoswDyUSGV17ZbDdz6jyS4GCu7SOzZir1Zbzd5nnh90
OlLfdPrw8uAOiFGGm4/LRPEKs9PMdYPPkfnCFlAtHeIeoQPRU/nmC0HfgtKzg1RmqMEKNDdorsyi
OPFBXS6ahyM0uQBV2TLDU9KA7a7N1htk8YNtnbZKfRoJ3xVga0G8lyGZB84AM6jOItdtGyP1Q1zl
SDt17gxg2JA6rW5ynLhlGeOVMnC45Y6saCi4izDEv+8NnTGVt8UShOgZGCCc/Qftm3qLpIBE06bH
LnDJW0T5EVEtRp4B82tzep5KsuNBKNbq4JHvWv1jB/G/LiYGrjL9Ze7CuWQivZdXK1MdOMKKpLeg
R0WTHxVgMKGYmiT61Vrv8sEYxRNTX0C6IXdNWIv3CpEtsynlF7wmOTOzinePm6nUDSxfltoXFJrd
5g52cX4uBAvw/jF5CNmWwz11YPNpiAvqG++lpH3p1Y92enF5XNabpfXtPhkTNAROA28BVx03sGS+
dSe9eTpBYN2jgTCRqh6/rV+bdhzlHgWfeAY48mqotRifUgO5OiIsrIHa++n5avVqpaTR/TYpVVnC
xv4cB6ln9BP0pDp4GE4Qj/Hk/gsdqQArOJJQ3+6R3cV6pGCbcKYN0h+AC+SBF54Zm0uNCPpQYS6g
p7l7EjZ86LK33/YcL1Zyf29HV7m5s6AFaNjUq0Wks4dCWJzqsMtRUJbbdq/vhFKU/KMwxZ3rqklB
lKNejxjT5gnLZZpouu3wuHIgVhT94gdkqsYb4WXCORDjW0nXYtKZxa4dIoD7PPFkBgulIhCoftJl
qlV3A7HOBWGnK8jGsSoHNfGT+Rg/oLiuFVyTTd1zksJmIgP8w/pn1BBjrQHHuvsLl7V+AuJUo7Av
PLaStbBu9pFBYWycjY+WAtA7GiyWTVxkIfV3llMBr94Yc/PTvhM/IH1+AJsONuDjCu14ovdCYia0
1R8y/Gds/TL4UBAT4oR6o14Br2/MDmPXC8ri4FDkLEkrSunmRvys0w332GB5dcGZXWlcl/CHLNNt
GlbWQVqeci+xZ967yBCsSt/Z9/iUMJGcO699T3lO1YqolN8qw/4K1bsIDo3O6lk4gn9548CsC1a/
DUI/vb3TOkntDY9gzySYDZePTB6i5w8WWzn6RbYD4S7rGH20Ve5U0xJid821bEafCOQOML9HWNHT
tYjje0U/cI4ZYGtIT6QyUwCzLsbJwWzft9tDr0YbbVTzZL2vE1NUGR+PNrtLk+e3Tiy+FqOShgOp
4fF22y3FX6vCnVvAfDVs/t4+INAgLzQbaz5rxehVqwjsSAPW5xfX6jqYOzmgq9zUq4D3eQNaPLuR
PVAA/KlYyahHsaYgcgno7XHJzY1WBnmWvNpKebuS6BE+HKI6lVTSGJnCxwive0+2XvXglyhU6Gcz
nzkxZeYfL+gjNazV0o45Zztbn9zR/AtGE8NHzP6v1sDFbh3VgzP5YN4jVqV6tyG2QGH6gqSR4S24
tSlfbeOs94lAgPxlIFCTxZTf5IKyJakh15VNjenUa29fou0ueZbCrouLeqja0QjvYYWjue3jcs48
CkHCROaBGfDXNOLh3z+4IPmc8ksVMd9azlJTn2+0LW5ZB/QIQ9IqoW9WbIwkkCeMF/A9ZuRAccgB
oEwFEjIWrlMRIXo/kwGj6aINI9DsFChXJKRqjjZwAKWdXueN7s0PND1m0LxjEVHUZezBF9whzREL
dZO2jHyk4wXz4s5w1yd8OOOVqfEn/QG+S4VMVik6TSdT9WuMW/cIk5kpVBgR4f1OetqqvuAy+NjN
M1TB5Ksrm3VP9/2tO7ybdCkZCWzhGhSQ7zdRl22Y6O3nBo2TtsLSVyiQdXQ2aZzHKEpBCBYyDoO4
S8f2faM78fmFAIiWhCc8dqfB1A8GZ1GoxvUskB4HPb9rSTIOXxLsGM/IDxakk9zBaI3swayEhydj
ygn2bFdXfcJ+Umc5Tdh/eXOV9/+OV3IL0sXOpeg/xz6PJzSGDAZrQsOAxRs0kqP2zSTTkH4jt9lT
QK7sMKzS4q+GNc+qg3hXFV42SO1eCZAQIP0SsCACxBjIJ1x/lO2IViS8S6TC35Q2m3BxtLe1tdQE
m1sCMWOluAbWwsXciyFoQvNpPhqPtCstzhH1CHji2pDm3sN+gv2+BCKbt6GhDRl3/DBTFyGEhNUi
PC/8nRNkSoFWoWVTg4Cfc1Ui85BFW4AAEEhdsbV42QONe+e/dhvTDPKVCXIziFDe2OegsDAF7j+M
AqRQBlGVRHpNmgpD3LfukxgCO4KKx6DNvBNYky1LhlapN0UDKDghbAicu/VQXxdyp/Gjm8ejtyXt
i35bbE++qgihTwoC/dK4LC08zGvU6/rWKGewR3TpQCY5uL6/nbqaMAXm16ZvrUhaOmG3l03pRFJd
wg0FmPuNx4H2DoWWNYgi2hWQPbdA3n2dMPqeLkg5UT4pEBTsOqhtLudD3Xma5okDgKh1qvVdWEfi
zHbAgFWwh3XKK5FzbZrWZtq4fU0I0Ody6IqxujrlZXDEvZ3H0uVx1DSx30x1UkWFNDjef/yGeMmp
95FuuWn3Oy66Gk0cNBspMtD3qgAJylDB0jBHeH4273yhCxGtzO+9+OK85rDXqqij8yFKy84T3PMw
XYJqb9XFgvUo9ziIfGvljXjKp6Gye5xYOkiu2FU75NK4lxGuu9IHKY5+3G60ynv4Pp1RR99+8iyR
oldqOEWXS2Nr4e6q6yIvmKBxAWDExbic1efmeQyMesIaWgPSp6lSrJo6ihK8xnN5RyS0UcBP+IHJ
Y5NvRhCDlL69vKlsDO34NVgEMneNeTwMf5Dkh5yGJfP69r84aGw52+4GtqE4/HpahClqdDygCE/E
sGa+BRTCWwU+aMutBnH9FbCsnJT6JBieAi1TtNFlTH1wxxqgO/EB7DHnxLrK9glcvJCsKFroPI9o
S5KSQDYWiLD1UjDNP/9Rn4rl4Vk0D+GMa9FPEBsweNKutcT0hwaFsQPkaHYq020C9ugqu1NdzGbf
oCnhTxoh8GsieTLbIZQIPWMihaKVvSps2iAKgQLUENBTdtLCOeesNINN1O0LdG+dSybLM2XkI2Zs
U1moleFsMXd5fxv7v7lub/k2bSEFfzepLcgx6nWfHisHd+3tBvJ42KlF+6RQRNsw2z6Oy+16Ij1d
lVsdCQOYqSiuUGAyZCeNJdht+vjLmh1A2d/f7ivNGCtRPBRF0k8k5VElqQ6Gl/kzmLzWSpJogv3s
/yCn189la8XXh3adfuiu6sissOLBv252PbSQXPTVccsm8te6ilJiV41DWweQoOdav3/qpI0+YCdK
NvmNL7tJhssGlYq1R0+hYpIUtW/YJQ0tM0H2ynstWFzq21hARYPayXX1JWBImkBMP0jwAbypsKMS
UAqe4oD0K6xvhJdSzyA/6REeC7bJhjv72g6Kzvs2hZ3iCNj9wPBc9hnxMDBbi0Ag6Xv12Yelh9nC
Hg77Uvs18owZoDi7yi2j7b1KfzRe70AeLrBYV9b6fwBvAOedL9W25bCUcrXi5HNeN+mq9W+kpO50
vzyop9e7htqdiE9Fvj2RYpSQPCvjX3IDsffG5gl2E+sHs/aO8zNruitJg6sjYqHalP9q2p5UUPIQ
DxHLOOg26taKNGZC0n03VvPdB2Izq0FS6YwLoiIy2PFN/yjVoUy+VTXwrXE6MqseLJTDtXqncGls
gEWP0aZOXueROWCO2YEzmPqvgrOVNQ1b+Gwvgeoe6Un3PZxBZvA63NTUEEAsqeim2uSjrQdzum3U
AR0UdZMtv9VyTLOEQm5gh/EAshvtdJ50FDuGKMMz3/4al3MiAn6l5iRzTQu7XWG7NwDs/4vJPHOn
htMtmou9f5wK7HmmjLogmhzvdXewmce+1xzAEB9mPf5E7uneQhcwZcseJwmeWNl3AvHCO2ImpRNz
/mi24F+h0ygAkI5byBsMHNEQ/vJz7oQZYn18MYpFiUk2BBFXqshxpfQoqKqHdnIYU3mdEi0cqOBx
7kPtuDO4yo3H8n8IB6k3Bj8Hlnz21TNviEVNLczylHqo1jGclRsP5X192vkjW2kfLewazskfdz1W
PLswpGGqv2XYMp5x/6Eam+IZgZ8hPYEmWqszBY4IAtPWME40fP9dMdwUZmsMS5fMEADioVw54Qyl
1iCyrVpoRSSoNRu5BU9N1LNtBUzWNAY2HWGcrKG5qBl1uhSnHXkbjfiykyZBgreXW+Hzot3KnKfb
AP3CHBqSilOzzW584mxKXba8Jv15PLA8r2uuE9nSfOmk57lIkA8zIoC2ZpeMihycr2rgyPzySKaJ
/UuFPaQb/hPSeloGIdNrojDdUEO9Ln+LegCjByYEi+k0LKE4oHpHEb61smNyMstJ6Z4x8B2nuaDf
MVa3Kz/oMnUlBAkqClfWXspgBdKPtye01XPZomTGXs/8g6OhcHeLsRAiXbyVaCfwz7iuH6Xhf79v
pbFrEfuUpA3SO6wXjgKAs0O+ypqrvj8kEIh54ZH7JlsjQvSbTgOka4X3ofV9yPY/wY8VWOvRuUKJ
HaJe6BJiZSqDoh9a0P5yzaUaM62lw0dDgeiE6R6a3wPdZABAyIkc3u0ZvMetm54s+qFbEdCdJjJl
utv+4a64rLdcp/QWPvbEGIJkTgKVPVXY41nZjo/GEWW32RDsakftVMdj1guLUdP2ul3wGoY9ABlv
FBq7iQd64cU3HQok0EXcoPRrbyA7xrVT1l0gEQuJ7Rj6qQNUeJPn/j7LzVPnEVfX8Tb4cXZrOo/1
Yv/xNMXijekRE2s1FGoOsg0EU4wD/upgqEhDY6IXemtrQaA1qAXm5rAPEGkk+KO3FXdWuiCkzQM0
UNBWttmW4ZGcbN2b/S5BY80Y5UmLVvmeRmARmpRVJUoNaAUP/vxHfrND+zzBZC7GGD38nM+YpYKe
wrPXsK8tJmjG8uGoEASfhbva5j7DoQI5dkCj9B2myXZ7ZcMJSgTBm2NW/K053GfPASP/E7OBxB+C
RAFmaMK4VwILvALzCxzxOIwlGqAk8c7Yhbzq0h1J6nyMfMjaz3Qi7tAcxraXIMzvzUs5q6URDjnE
hRXgQwjURVfq4Epk9zftDRU+bSiJecw98WWviALr2mdyPs0K/OXuV8qBwLvFRLsail1SvqMO6KAF
xyf9LdNvrzwMLQjDrw9TKwigPwjbeQOy8mnTSa7KLfS/lmrq/iQUNKVxxYLHecw0C2RhVI+Xd10n
1vRxsakR8a6yWdT+gpht89xcC7sS75a368KhqeAORy8laAcjuYizY+p8ipvbF3/D3T8V6Mmk7CBw
JLuVh8mFehovoMd6Pur8wYBeBo7nqFi97W3eLjv1GX8utbP684vjmELOCerwoK9G7ONp9uAJgdIp
3KnY5gr0H3J0km6DmVlSaLuM5NDjLC9IIxBGgLVg6c3p9XEfBVxHQApfV6Rtm5Boz4tK4Upt8cw9
2/e12uWNM49IM8AuzQsclOTqeU4sc1wf7kACX9OUlE+TjR9UY0CBeZGLxprAfBVO81m9reo1UFxO
0VvR1C0O/jb6/ID9pFJfeTTQguYat1aBtD5yqVwfer2Nh/wRW+9NTGSpb5u888gPyHwJyVJYnhWr
GOM1hZjJdjjEK30RsaAOAMEM37KXk0xrM6huLeO8GfDvOzICSWR/3RC5zWk2JZE/GY9PpHU8sX43
gJdkJZ32EU+mOkxGjYGElUWwZNMUqBhEUIkWBsQ10WwBxkoYJDFwKbfFPm91VEHuSC/UgS0pYIL1
HRlWxxUteJyygMXik0VXN7X+5Vhlf3fe+kcr4mx6t62s8jLG/6Bb0+c6guvak+2l/iQBKovlbofb
Jy8t76mkmm24xiC1eQXhi2fpr/cqBg5ff801rE4CO8OlEbZGRhXtp7T30Tl9mAtnN9/oXaTHEtDm
E2gjpZnZf2LJK9f1Vu3V0LM9HiUNXGIWzRkjsPTyzi8t5JWiFHCBSATghaz8HAqpo5vSXjDSql7l
J/ohmOKqtsIxATfMtTAWvUZweZA23UowSh8jKOEEpl/sSznnQAOmpGouvVqZQYMU+ohF0Mpop5Qw
A/KQF+uJqTEU5GW6JII+LYZc7q4vBCIUPQ+TXWqeN6EtzXPWZM0UCnOujELSJT8jxUM6NZbZ/MgK
nzQ7j35ImeTxr1y2ymrh1XYdTc1VVQrE+maBh/qTmegd2eBw6V6dhIDH9/QfTocIYYbLdy8J33cT
JxVPaV+fRirsxh0MEHTAakv+qNAxuYnnoP44tvp6JSFRDnAPCI6sJ4yYc0mw/QE1lNpxlEhHTE+K
d4WxzVtJf7h/VSSG70Zrw+v4iaSLsG0OaBT0rGFTVD+KuF98YlSmQoK9g5oG/YMOvOjgocCPTuYK
bqKmuZ7gdSEe5Mba1XS3qL9cr9UH4cZE3Api9gmzn8w/AaTT+fQ8GQTHSXL7jf1wNBm89BYTN38q
a4EVkmwNKIyGEWsnlba7oDvkeDXCwYSpPa/cRlrytXhUCXHGsgNFXM0YeiP97g/qm0670xASWOrN
dswUiukz8AoQK5821h10nNSF70pc7lR7nolEv+HvecyX1dpFCyPKPLIubEGbkEsyuOg6UGTMYRQL
JMTvqPjUBartCbU12x/KwBTNVy6P74xdvlbyxRfnIOF/ht1Zd7R+pyCvWyFyFVWxBcGTROWjkcTK
IGrgj8Qdb1EVTHoaaGMdM1PFcpdYlOdLIQXoyJzh/My8YkqvVYKJ07p93JXWSpDPexjqlWASg8u1
Lii/t7bu5790XcuyHJvj4whgCX27R84DampI5cyEGKpysegXeIG94WJ18e5Vw1isFLygH4I1VSPh
umm+rXG3Ig+x8fHf7xYWX2A9ltCDppaiEOPjMe3hyX3UYCF3X0PBspK6TjJv6p+oM81ST7ETHExY
pc4+wk/m8GPy3mIUF5lR7c62XGpcOnoclgGOpcR2Q25p0+gqAODM2Taw3D809Di/JQQ4DWL/ucsY
ewDY2njAD7w220ooTlABTJjTUjikBsZrYaH87XtMHuJpfzLFWnw5gF+0lyrz8bHWOoYriibdYA11
w36a/dXNBc6Nswrlkl4WliuXy+LC7/S7779albah7NqI3Sgph6MFd6tlPxhLGQVvaDTywut6YEqq
gK6mw+lKf56zOgC9GEbpBc/PiDS1/EkJRoZzDTQyXcQRvU33Tr2Hz2eCvPnvMjLeOlm8tHhMz/CN
g4TFHY4HAJdLryzxo79mP1V4sZGMces33qftNdfQ+eZTZbqXKw/1mFFvK86ggXO7hoD3e3GELcY2
RPdckckL2Bsusg3mwEaV4MF0NkfGd0LcVjmzAVGvu/O5HM1vNTAfEHkGgMdor0NnemXfaQPU7fmo
7Eq8UDAXjqFk2K61mfOJpe2S3BRDibS03A9BykZuvab/AgscrQWuQpbusqBMGa/d9HObZ0SZdgVT
AjSBOvKA3lJNEziW0Wmt+lNW5zr6YUMS+NouhQc6HPaD7jCQEBb4vb/tJBi5b1iRdxkp3q0P3upE
JXPeb8rMBT1yyr5Xf2Pz1U55kN5Te6rIJ/aQ64/zj8Ds3ESblJ0Fj5NfD0sPtRmJt3rwFgV5YoU3
te5eK2KqkF7D6z+kEX3o3CPcQrjWMCse7CcLEADppFEThPPnZjczbaaISWzPWCLYOaMQ97l5xMgj
rfjcMmRPmty9Ww4Rleq+XvMwoBa1l1qNBK3/SdJ3ECys5dI5/IDPTJjf18M075CsLtPNzvnDG1XI
q0of0BRD/9ciTU+kQZrF7E9Pctrpotco71LVakUesBJ0WLRyWynol7U86RnjDherHz1QkQJqkiOT
IsByPxOGB4Gxf6/oeFaiOMNpq+R5Yvw0OM6qP6PJabPjAMd/XbNSpppyHaUK03LAhLJg/1xnxpQn
SNXi8SnkWdGNws1UsGGmu4PSoRChqde4MNkh/ZQkFMWaVDwY30a60aZCuv0ODlXfqV07wpKQB4Xr
MPlhQZA9NvztUmAFULX2HCCz9j4bPSYySLwHM7xy223T7y8ahC/gmNadVf7TTJRdfd2EDzdDjw6u
egwOupY/I6/sbgfzqx83oJw0mzX1m/g8n4W8CXxOijOpHSEobO6NSffEaCjim5ZCnBvqqj+MsJI1
TngOJ7qf6UXqPE0Hu81s9Yk0PwrvWbB4Zew/i9pis9L5AXKAQEPqfMaCEJCbZ7XJDjwudwfW+gzF
3vMtrHuLmYfaT3IL4PVx65jpWvY0cao8LJcu69BoxzdhXWLgSwxmsdv5x87+lYLn9PahUdgO625a
09jT6Fczloi2SPEev1re0kiOt4yXBDAGMDYnjsgDksIvpaxrJ8nGQ3BdbESqX6j9Zs2pMC+DvSu6
l+6dcTnIQfkxM3twpd311rN44GZP7Tsfttxzm8qKu4TQJUHxDtpvX87gtmA1Tf8pwYPVZhOzIr7m
k6hjvyo5ejinGTIkEGU2BvUK6ezIl0llEtLXq9bliUEHuj89FJanBH7+UlWfE6mT3z58Tx9ng1+7
GjPPoT4yQdEbBC7MN6AqIEa40cyTTIxmCkIY3RatPb9arkDLdlNeLUrf1Syip/JV0NlnKFIqU76x
r94B20Kk0/Djux4RhD4Qz/RKq1VsGC7hekU9KU2XlpHGTUR7Vp6Wq+nzsj58mo8G75GeqYFn/8/k
Cf57HzdQ/nlm0MlYkvGP5p9Szer8knFQJ/EG7q6GfHpdPkTsRkdHb/koVjf98Oo2DM8NYVk1Ypzo
t7SfliLzLDXcYLJt/B7ynZeX3c8StJmaUxgOVZYrQCM9G/oLjjp2X7W9BzvKtq6npl7tk7EIzcmj
jlsua/sM9nDzklRT2KPlsq7VF+CM6xoVqntOn+7cetdDTSfqn1L6A47q0azCgDcPZI2hAu5gP7kv
8xAkV0l5yv4kJquLad3qXpjZh68R71HOFPIlfgE1FPpaxCw2vhjTTL5ZoJmUYhjYIa6KbgOXFD3F
RZvxGn2lLjz60SMluzubYTLkKJrVSpRzfQUtoB2o/jARBU5HOaBoRZJ0PhQLxx+fGmv6BBqh4xlS
omhTchysWNAMG+5jp9UYuVJxTkkQlmsAWujg8IFK7ZaSfZxY/6n6PUhO/pXaNhS3sPdOS/fX/aaq
lwfztQ11NGSEcG6P7uGTBu7Q8HTgaaavbz3ill3etUhVcBLOTNa7JeQn1/VHB5nUkUXabe4n2OVN
RnU2cia/SDVL6qYIcSJHgc5buMdi77K4FAfWORnf8SQ21FAz177v8c23EafyXP9UmFzydmezyJmJ
+RbrTC4GNkq2mhCr2d4JPTvBQC4PsIYr2L8/T1rHAeQiQj8JPYY8pE2yQj1tFn32K71wV+w/ytIs
hujDFGy4YDI2VKiKdVSxKlshJNxdrc190riPzlP+Y7p9MP2KTeBSXZpSMnuKDEhhm7JE6oSJ8TD4
BjXPLF5MtCgVBGEOkE++AG6fv8M+YR/29uCfOmPP6HWkc7pDUSEF9nbnTO99OabUAlL29GE9rrfg
SjC4EkooasMG/fuaX59NvKMc+w45SuQHSFp8oFscoBx941I589BdXUKyXVsWKRxVdPuDQ+CtAG4c
9UNDMWHEnSO+6EMFXQyVYs/3MOAdcQ/7KguHHQ94wMPv6RKGo7sRgkdCyPLEQKBF5NHr0m4IE0us
0ZNt0ajL3ubyGjIb3iDprKho4r4YsaZSa5dztoYtpJRIHxZMX1NxWxmcYafcLZFI1e7eu9KtKzYV
6fGW3azhGCaOn4bjsak8tY9YVBRb0Fj1ZykSQeqDKCXPB/2I0Gub45rTyOkkp13yQJVljjfqnlJX
+v8rCUmNIbzxJ9eSS+qr+2ZJJ2fxRTQyHoo3miwGljN7td5Jx0bs000+jOaEL0jtp15l0yAlkE9S
r/W2P6AiSGp6c0ttJh1kCrBIrtkBmnNCcn4K2ISdU7kDWtxN4hYb0j8Y7OfotxAc5K28IorHGnTP
f4DnOXjgawzFOh1i4yc3c/0MXVIQ6XK1byTzpNYvEt2gxCAI0yoHPtzlcT+RkxSu5Gmu8vL6gtGj
N4DyMnbqVdu7/MNYlucJonn1lFY9Ty+HGjBsOxQVmOal/klMvBUdsVnJ7wknYlf04/L+FHL++9rC
ERZtHASDYeOD0pKKgWztr0Zdv0/aBjxQJrlbSfavuDA0fgQ7II1FNt0SdwLISov/dYBuMb6q4CSI
FXSc7MC66oMmqHhWA7WAnccL0V6vmd7Bq038jon4lbaOjmeRljB8pCrOfIczu+ouu5rIjjkNBwdl
qclc4tTOFtECl+YYtEChUIZ+MxfHClKaV0pkT8e6NNzubbLLPOtzGETQr5elvqksGV2BFJ3cZPVy
CvXBpMAzk6T3n/EzR4OJr0HLqS2PSVpOaxjeS0b/4wz0i9OvfpMqIWN0CQsE12V4HfoBTZ2NUswm
dDgZPIlAuDRYzV+SS8xN2WMf420O0R9hBwCfi0qwIPyUmEzrGeqRBOsCPlfbdHlLPdbvZ44H9qgA
iyUQ8SNHR+D3SvjVV+bFTArjfar9Iw1fnIXsAdTNNJd2RVLVDZAX4r4g1Uk7duORHC+Ggi3Nnxlr
X5B4OSV+m3Nu4O/qUqzit0BvzA80AqdrFD+zPjxWU2LGfQS05iYnphN3vgGeCAZoU+zsw0DAL3Xc
DdvD57G3TNSQ9AgwVSbP/frNo51ZYhaxn7GgGkFXsaG509Dhq5jOaC9LIwk3FKr/R82TlhtLWOle
82ceIKo2GASNTIivNTEZeqe2qMQIWfLvgJ/lXqP2Wx7++TH4iwI8gA20zJMoYGy5SVRHXHN83pbw
D4eCdgdc/ILn8MD/GfijjEMh4ty0jKGIbQ6kIYpGg9OkD2+t/hRtHANBzdMW40G5w7fylphre+BZ
LbHRY3RWLq80Yyjl+HAqlecE3ChDVxcmcDVwQQtxt2Z/eHWUQbaE1GYk/issAKidmpQwMeTaNR7N
8Lzl+oL4IdVcnliDZFdT2Lj+i4/2P8Qw2+WlLyJ3QnmCGQoxQFnQaIav88sHUYE1tLnqM7A6cERh
XoFIF5B9au4TlllwJlXy++i9IblvCmwV5O8K6CraarBVIOOfK9kmrqEM3husdVD9ZN1r1v+Z/Vu0
ZqZD1TlA6jo8Te1u5Sx6uHrv9gjDwCprOBwSjumeQp8yP4I7D3SkZ09COGLABoAsc0CUIi4bjGPD
1AcUqSyuWyKhpXUaGPwtjGkBliVn+Zjj4CplFos3P+3hUUUTXC6N9pejvyPEkSzx5yYJDPqqtnCv
FBqDgLvXrrGA+vbTA29TyIVrzHjArVH8LF5u8FY6On7OfDFJZYImRZQNfdD1HmlVBdzeUiG5lAEA
LoI/WMgaAAkELu74447nS44Co2OF6/AGYKnVAU5US3y4hhgN/WVNQf/jk+/wrDYNauOxcMhmK4rr
jmR2QIg5/QQVzpp+fe57sky3JfVHSI+LHWrBESQF+pwB35xbc2M0C2nJdYpzgNdCVSRlMX3CWdEx
dgfOKxqBCUo/nxG34Px3mx6IiGEhkh+779yM72rpeJeM5JTxvUyD0JeS15k6iOVTN4sHMnmBhTFM
KMpKYI+uSvTViE4f9O/TLJzx1Ll683BJu08l2v3RVvx73/I2eJdX/Q3wJfNJ4DJ6UXlIq6Dy0gwR
S/xyc2g91lkZgd0X7voUTmEbSzSfENEbA67sO3PZynpJV/FyJLXBmgmIhJggCTQ0X1r+KU32X9l4
HdvqYIMxtOoSVuO6xZbnPi/XFZ+2lVj2cWZhezCbTDfu/z6elrBnCQSENyS1rTjy2a/4uzoM21x4
UvYv8KvWtcRzrCD6Xv5Bo9nsQ0dr1eWXNaLmEIKfZRV7btTL9tNLdDQt8UijWihsP230vYFAbCne
vwxYaCLU0YzG+hVHb5DfxgONITa4enaMinD0aCE7YLEYzimJtGuFC25UW/TGOrT6vqsfhAoOs+F8
EfYXgSU0hcXxmvx3nZ7yLcRUQGcgwghDYZUpyitXsc4D8wQRMiLf2BWJIIKTFGxbEFzDWoProty+
63fUA9Ve7CugMlKzBJnr+pKNJVQm5dgoxGx1jmH8j8A4on/a9VJFa+cGbagImGjDRZyFCrz8/RKL
sb2vYZN+r29PZlK6pmMkMma5idLBIlgxFpaU6juFqXtt2Y4ukUa8DGEcus9UqhpNG/fjagmOU0PC
BYrOLn7r/g12m9/fNcLIchNsABQObTbjkBOF1hGgsWafOA21pfUY4DNwuDOts1VcHKYOZmOXwk+E
jcHL881KkFUfnKD9NjwZj36GHnidf8usBJMsA+9nGichm0s5sOJTEarAJH6ANyhlCLqGyPeCYpSp
I9+/uHucgrb1MKxrtQzXUGrubWq+AqEJj1poeWXL0kt+LRy8al6JF4cFnW255CNTsbOk81rGK2N4
V4Su+Xo3yhcOOUJUZPR6P2+fePAn+ZqKX/wxQoQvDzPQipDRDTu8SPGV4MZT+JkHrDSo5X3kSCQx
EzckKcH9tnUAyZFw5lDZmZgC1xb5h62Hslm58+U4VJoaVRhNUSNzxIIjpuRGTC8INsHveA7Jgmyt
oW0RLif8eCsNEwlQxH1l1bMdA6QPSfW/Trt7XRkJADLI13XfdgWuoeMV53Rc9+DCOBcJlit0FAOK
JO5K9wcCZEph3/QMWBWpTS5F6Udhau1duwYEcvUDfR3clh8qSkho8O3F8HteUknTtJTUhYObn/GW
bJ+eKON1ypDVKvBy6dnWk9ko/ZaQe8aZKL/c6F1zTQSyVlcOO4d9p2ZKej+7nB4CX+DYMPASLckB
XAF7ccD8mh5fpPbXJvAaba2KZFj1bItPHfsN2Szqx/RtLtEZLjsKXVTejEgg6Ize/acNnRtiTC4p
zqc44lQMWjQ68Wzro/rn1rbOcrZ3lxLn9iMqa+a7nCPcO6oBTOYHQTnFjMmUaOlX5LfHkcGSlIaJ
UT50lRtJayY5+7y9LS7Yi333volRZ1JNgO7pOwBpqc0uf9Tsn9P2uq4MCdL6CeWg1A3ypL8j0p68
q5HrmxXPDw9AWCFPvJ20MINdbuDo+l03DpWfQEWtCTwXs6d7AGb2K4Wu7tmwp1lNuX2GiKiUO8eY
oUIgdPNhq9GGsfxtbZvHTrhikubDAFCqbiGejsMCdSfoy8anAkMEnBUJj/61aJ50s5/MzNDW3TAL
sHPpCPKHYTnQKuKykkduJ5U0X8ifYQ0m2dpC68yi7ZCMt1QXpXXBc+AgpeJ1MvCWs3JHWhrpVW/l
5mJd1MKMCfpeUg5GPIN9V6ptg5sS8vCmgM7QIeuTGfYzSAA16970qaNOCqPpIFuNmpfhRWveZz3W
6akxMvUd2E3o8YWKw/0s74cPgh2HSgDVEPVD/9fLqFnEkYxY1R8xbdOj5wtUMxgGXXqUV8/0B4aZ
PX8aEl7LozMZZueOxvY995pBbugLFFTdFbUGvJ0mzl4NWdc2KdZkNxNC5PAOaSHHdXNMeqIIImzM
u3HOyHq7Oi7qBmbH2jS5xAi1VJ2nW4kQbQyEleGZRaWiaSQwR2nsX+E1ZkVMYwEsk4cRy51Gg/44
dxvPYy5++yvt7sdwchCBUmZjCssnAvf2bsmAmGfh7/S8L6jLcbSnPsqmpKLYouu5hdLjqrYOAB4/
R6/kXceoBrKhw3JybbYhQqG+OQRGsUho4sSbBQmz/kWxECtDlYKtoOP7ohHAMf+sWJPAsJfY/Vdb
5Cd9ID8mRuAK8RAejtB65PYjajFFNH6nFIBrJrFOCl4pBE8xLxKTSCPqaah0OE6CEYby7t86vPVz
C/T0NItQsLW7XK0CNunfQeai1LHtTAQmAaXdJKzZIyWWNC/2c9cbsWV4Cjq1bawijn/Dx4yQDofn
H9PwZyC6QDo6C/UvlNxaEvGSdOejKHvTOB+kWKi0VbzL1s6NjDdFWnV8Mt25AxMGBfdRQvCQfwZ6
sYHSuqBKz78MxJR8XdPp/P4zZzc3R7moR9FzXQPLbnwpEemMJCEj7V+I+hZIHL85u2WV5m0X1VLI
GQ+4s193orL+bRxes123Itlx084TGMxS7+CN4gWYKtwzUU+J/A1Cl4R2stpK8fxvnjxhFOBxO5YR
mESY3rzlWFoewQAZP6mEvSEz7W9UsqIqmqJC41hFYIncVx0YOPGLYEr5DszI4j+7ZqPwFMsTLZkT
7n9pP4W3PGPCDf5HCXs6nuKE8Zukgw3Ah/+fB8lcpy3m6CYiyUhqBZfDN0B2cizlt7YHCr8PU++I
zdqm5zQBvFmP9jpjkATfytCGfQB5GQG8P0BuWr/9R16quNuxCyTisy4gveVHhxDc1C+P0hQBi7AB
rCzs5dZn3CA2L4KjxtesJjyqOxGHVtSWfwmNdf32O4u+W8AyHlVXjoQ1MKq5gOzI08ijQSaGOLg3
PCj3tua1tEtGJ9qDFDDu+BlYXwObv+mmUdic8K0mIeyf27t9vugQ9az6pRKy9F6EJh8rhqj1JFcS
ED9XDkvI2uRVJwcQRmGuUUsX9iaAcYfnt8IQgLupHZgJHssYjnNEV76DL2T+k8IbkaZ7MQzMCzf7
Bpo6VPHqf2NK72k3YVgW6b/V1gMrUPjg8jpBXRdhWDYAy+w1RtyQmvSvI0o5XNXEdC/hV9wUuOJY
0FFIM2cxUNqGulqbV9vCAimP93GbVn7xIWfXBmR8qIXoBCU+wyAQ0Ko0e/3nKTaFhDtl5xHrMsKG
jUFyppZcaFORsO3B40YK4MPJGa3u6BsBAezx09apALLS/iyKikAAdJXSvmfPFJylruWWtQ0z+lnn
iFaily3IoszO+QynpwN0P5kSOW7YesKtYH/lQqbwmHPVXZ0CBp4WHZ9qjOdmhN+34dnqft3fPQ0Y
8fhCmASyul+fN6nNqXt5EBGxFZG24ooxHMV04gRpqxFMxE3apE5DyY4aOTqynuibvhPlYynQ7FCO
u1OFJDZ17FXZKIqmLyGRlgL0xfJu28V6l8Dh3pkkRh9cGrRwLs3bfqDXF5rdxQW48eHCbvaQLeuY
iaX25xaxpx5joMKkX5iKbs2gLCsOH3fQ085JWJmAwtz6P7J4fr45cVIPH43wt/NcaigmQTnLDOtA
h0JGd2SY+z0+6ggwKf2TYRa8x52S7+cpb94hvzAaFQCQ4z0AbfSU/U3KOeY4vFSio1+FASiXa53B
e4Co305Cg80J18jIekmle/qs5iRc1R7qViygYxGycqHeuKvhZrZJt1kY51e2FIQpXrbDeoKwmci9
xen+1ACutYaq/ynH/51dZewN1NZLrQ9u0BSQBljVG/b9JCKQhwmCZAoFVpYeEQMdPx6Ejmzrep3n
cs4A14Vv7EDdH3R1aU8Qgy6nfFSzyQiS1YgsuAzq6RZ4qgcO0UKRCBL936YoA7xu2vSBIGI3Hke3
WLxXwZ72DxbdCloZtydCaieJgrAlH8UuMcjm0vG7nXmQiSmXbzVL+Rk/cYWNtVqsGwCjP3vIum7t
lJpp/sgZrfApArAoftGpSU3464TlUIyQmUWBJt7flHquAxUO7nA92dBOHeacMBaw5CYzB40ftudZ
YqYnQ5eL21d6RtX34cEFH/X+XBy+yIXMH0F1OZ/BI/C5JVjENOc8N4Fg4tbngLXsqci9/ywDwOg/
QJMcRPutOnPnw26BktAaaPMGOzidlyYrS8q14jbro+PspbxyGQbaeHJOk4iURzusWaGkFH66cEni
NjaNykd//wweS4pMDzlbVG7buOZMiSvVEk0FT7uZLaTxxKkdOuAhGF/vhMGjvmExbRZFmrN0yMQC
yMXcs/4fHLwWV987QPfIp6pSOyi/iVnQcDoXyeWYFsAWI+bRk6V3NCpA+G1aGpy2k7YRt7zlEGtL
RYEdz44MZHe5ZATf8yTn/Zecd5Tcen8Z0XNoitu51A4ll/ODkb69QYjROzEKRPPvZawaNjJs4maz
WSt4HAKem5EErtobvxUXJ1HplOr9rqQZax+RoxZ9EjJ5sXxaysiyIWcnIk9UI4CJDSR8DLkmlXik
XdtJ5PeON/ZO2zjR1J2QtKmuW3QooBegVoFrMtn1c8q9E8BI/QAJjGF4gOJC9/U7poFuU8Lu61GJ
r7qB7/TsMTtUDYcm3j9Fs7mYleZ+sajhmnI4j9zu/tBhLHGWc4labx9UpQsZO0Vs9yr0LUgl7Bn9
7lnsHwp0wGklWDAgZdMUK6qGarOT3ZUMlV8e9Dm9yw7YYakU3zTDQ8e3iuqueati6VqpOuB8NMw4
R79ZBOMXmUEhI5Af6ss7rhQNpcCtXWswFODO2d4hyzb9asyntEWzWBxj/5kMH3JQjmgQ/bf4Msse
legbOoSDjJtXYMDHb/UhT/R7Htn04ilzWrhORlmHtE4N03ZnlhUeBoAJIFA+r/1WP1vuBZEXFb1L
wuUV44LTKI5AT44J8tgMYe+q5lM04kvT2l/g0cbYBa3e3YPMHAzrvpO8o3V+NZ37smdsTnw5eF1n
qoKKSDNIHA500sxf9Ogdpvt9EBl4tlygGlvLEvRi6bAxetaRA22K0wm7GbMya9MIo1Jrc20BFC5L
0Wqx0uZqCeG8zWneuLqKPJA7ZJC1I/NivRnuRWRJrib1uVy+BTN9sefBfe7/EkzOsa8TZXPn1RYg
RGiT4LuIviJudtggxlDoD91kS4RST/PGo70gDY4F9LNjYlv4nqxH1YNod3g+jyTx4NVLC+IspN3M
jq4iBZdZHFwidwa1njIckIKnz5Ck2eqHKGvjntNc+mUruW0SS7kOHA9/q4YDObFRjb09en4h01Kx
p/j5QoPamC76iDMk8VSpeIcVvh4aJVnZzb4lGFGH4IrPsHtfD7CKeFUV3cEVWI1FXwoOC3c2AKiG
X43iwj1NGhdXGdKXMoWvhehs0y5jtYgas3Y3DHtCTBUZYrkyy2uC0c26iSAiX3UV60WWctLWxMxV
aLGcEv3t1c+4dnXDrETNOBtVIgpwOTfQ5Hdn8oitkWy7ivc3dhvQMc4ay0XVABvPPX4Vt/U7m32o
R5e4eJf+31sU3w+8Hvg926nJ6BbKBdT0ZzyEnu7YfaYuNA8TNvoTiRioDh90EkJveFQxtyf9DJwt
du0qt54trTA+PYM9Dqfrttv5B8tSFxVIK21j1TPklhHvMa1vJs6hlNyuUW7yCmyxBGGbtlJUFUEk
3KdpH6THGJENHhxH09pxmy6ZTaQaZaPuEA2uUeT8O7xH0ntfvaZhT6XewJaNEVZv9YHteqFyxllq
h6/2urhRrv5vcYZjENLQEkpDfOrPGkYAuNpkbXr7BYHnewt4/Q/PeC3JXsAuf3/eCzY23XEszlyj
BCiXFogkEVBfhwg7rcMfel/fxo/Bf8Teb1kNpjftdPf+Ue75lljLRhc2ZpvK3O+knW9FJ/69ClZ8
+doe7qmx3/8eHxDXF9jdYfIakWwCGLx3ETqwSPin8solBTKCgCmzUbsLLobV+e+s/ZzaFYxZ4KnY
uXe/4Tz7pQRC34oUzKbWy2TClW1pkiO6BLss0EzNMUcXUjTFlcHK0yRlDLhUL6Uk0lCqg5u0oc0A
CknognysxDPoLi2pjjIakL1qzl76vcqU+cBfdixidMlxu0kA5RpfDB2rsghiiPU84PwgK34Zqp8K
YHKkvZ90QRhBIQfgcJrUnn0wyhvSPrlwHRtiXP94whwfacxw4TqDK4i+r6niSdwoa3sCriunsr1K
iDSutr+mecVrO6vQObyKq2ESP1xsIofjEF8K3yolbpUr2OiP5QqFkVE7t46nHPfEubg1iOyB3auI
pDb8w/5qu4rAYYmGYOFwb/BflFdwchz/S0GUzHGvf8ZBaRv0BA+g47MiWfw8gPp+2e2fe1+7qHV+
gOihhHP81hGRLPI2OP2RRBp4mqb5QlFKA3lwDxkflgm8ErYhU6UhSCoyj2qe19pKWSMkpgLcs5yG
Wz9teBLMWsI8quGGOaKyXCwhQaHKyA6yWLEwzCspN6RmNF23ywtUBoVJr71DSXJRgLrHnmAZehu5
rD3zbJ87SMsBWbyW2laDGRvXBu1dXlCLmgaFTjhKvzIWOW+NGbsjOxQ+elwIsd+aOb7PnNU5aeNC
5gZf4gGNflP3IQa/bM2I4V2z8py3Gvp0+m4X0AQ06XuPec/0710d2+Q0j6vNDHf1MZn2Tg+jJi1e
X21XUx8R4v8UiqWuxjzD9EK2rE+cY46/GsbHcWITlt5Pxx06Au8g506FJhLHUdq8V1Ldsst+wP/J
qUUH5D7E+6D9b5RmRA9N01JWJTdgEBS2kydw9NvMvnoWPz1rncPUL6uDNfOWNqhQJ5wX0UhVlz1n
NbUVK1n8+Kvg3TojiIQ4p6tCeZ3XrG5lKgyc6ZVcdNd64vgXG4AfdlulHCTBdgpW3DgBvVNgydaU
lAC8JJAOYZVbtecX2E/S97JJdoO21BC1zKezyghhCSQTTZwxEbDyo1xkrIhdtasLhqr0mXD2PII3
k8e5Ap8Jl92x2Qc2c4Mv1ozEF8RXK4Z2YGh3GjfzU4klO8Lkzk4OQ76XJYFbcizcIgWslpY60ah1
WunX9ogYq+WH9wFmwjCzatsaPigR9AqOUDyu0ptAOPaad3p8q9kTCjp98FT8FnFt3tZltvIEM86K
UlxpORFBk/OwFSKET3ICKkSSkmg/YikFKrHI2dyja5r4ouSCEiiv6tiwzg9BPi5KS/ngG8GoGtsP
muZxHFuZCVxOP//Mu9/4yMz6aO+yXviFX88otgDQ3lP17oW/PqJPfEQ+onba1MaAnFD096wONLTQ
UbC7OmoFYdECFuy4A6Qm97xrpLJ201jhHBj5sjAaiIZosmG2HQFV2mrHsUm3pG6ny8IwPAJuR6bS
9jSCo9ByhrRvxyLqsj8/4y356piP8AArKeYyn2wHFf6mnMO1y1JHhk2VkPtDfbJ0K2mopWptz5vC
mXJ0tN3z4AENBXjFrxvZBLzbbsmwvJm7ummlIMhfSs8idfB+yHs2+BAOCNxnGmKBoPtDEUaXaDJU
rYz5HPc9IPOifRraR2rYShn8uhcHq7Fr8vwKYzrVnabPAAgiZjVbD5zEioHtCvkzmg6ejWMo2AUQ
h2lv2IG2B3f3NheKnxYoCcCAVEAxrDrYnWhjK8nkgwuH9gTv1PXP8BaMY1DwbNSvaFl+8BJmREfu
bLvHGsIZF3zgdEXRMHHiIfF+zj2J+v07aROs/LF+p+Zi5schUsTE/laRu5S4fxB60Kr6wepemQQG
IRMcS8KihPaxzoPJXh6KiC4ldsqVasXqehiY9FeSHIa928StdbrX0WzVG7QnU2GepVaGvwMWrxgX
b8ixDdAG3yUWTNCSEQaWfpOwXNaZ5HL1dU0dAoW3ynREoM2Zey9jHi5y9WY3VFlSfBnxmmEMbB7j
8UPFF6m2dyrOCiE+YnI10gtHovCyYtFG/v08W5syLJaulDzIxVd3KgRyaVVwr2GGSvQzGxi5otzt
C93KLeE0emHA+1FbdVY0WKVn5rsbzk0EVesIUyEtKTZRHJZHxKE/p3bBqqvMYWzjUReUl1BjDQKH
4030UMa6fUdZnRGcB3RDVsuGFRbWk98EPSzTxn+lkjaAScJwHa7adpie6JIIWilqxDS9F5Cd3d1o
gijTf1YwjUT6tE9fn1sJWLoGKp24gNt0FZ76NxdDvnSMSOtv+aNqHEDqYx4gMSkrrnqpW44eS0jR
tA0xV/81EwDT/n3P9cypotNh/Js6IBi+sjbLyWdVT3zEIDOLO2OuiOJK3S464xsBbjjI2FeLouIt
HyzBjmL2wscNnxsrwE28md7qKqzbMsSCg3vEatl/PmWf7DQgXrqoPx4wcBOzKOSyuYWhomnyvBTS
MIFpIzlVjjxRi8izBwuf30SL0SMf31cd9uIIzus7tIHpk7GdtNZ8rZCMgg/z+Y8ISLTUY0CQTj++
SR7zbDlrs8ZrWc/biy65LXgLlAQAy/IwOJDZjOSmK5Ci214M/GMTo3gOw0sNCSRwRR7B6jnQGpRU
8LR86PEu8C89sdtUIEBEmuVJPN3ncaEMLSUuVn4ZXZ1Oz3+Yzr/UrkTn77zocizVrvWV/OP3Njgi
r/gn2qLZB9pdJqIkcohcqDx3Y9Pb97lhwvW3RoI2ktwcHei6pd6htAHtMoczpwv/WztCscq4X8n/
6frG+eMUHjJkyLwV61FmGZZliSBPUuKbSNsnKdPUIMl3FVr1CcGRu53m20IJCP6n8Bvfesks2za1
hNRh3kY5/adO8b4lcsgUhb2I6AWwTmvcrJrur7p/4C1dg36j+PK6OSo4hf9XKBUQW57g8Q0S/RHN
mE2Q37xGvprcaT+TGKsG7Vl0TiMJFo1e41kHfsEu9XtBRuRCTIN4zOSdaXJ16ERTqbv5IuYWs4BY
gDQjk6ZMW0RhS4ZvHyUo5F4GccFNbuhGoamSpM6Z210cI15udSjBUR48M+kaCw8GhEreWEkD+EHM
pXWx+ppjT59jB5ePcjgkmRc6mqRTIYpudAzkpAUjCScy5sOwG8eRmKsBqug9GQfUHMWEBV6l0rF3
UNJpaIR65DlVxSYH90hUoyPPDycenxSsKUcr3SHGKydSi19mjp5Nlk4Wa874HGNeq9SvPuhrFKjH
nv7MpG4pCbJ0nX/OegE/QeiO67QRg8b/9hxSHgZxXIrghHP/qOAjcDTaDfaKfFUz8pTVMri8cZzD
1EBil+DydI9yZfyTDpTLvwhbSseIxQucZSc9/fZI1aLDvl8+D5LE/SX+0Gtkw012nvbAmkIyGmOT
dJwXLw6EveymXe8RDNmRuy4SBVUXcagt6+QrhWGA/WxcRpl5pBTCZFN1nsihenfORtAWDCI2Jjpg
6lAOkEOVsYEUh3L4ge5MF6gAzc0/QW/NE2kQSubl25wWcg5fdxibZYgoTep52mWOfYh+vcVRKt8v
i7aDfafGmIX1wgGyNN9X1OFr9cr7HUr4bw66gfk2cul2HuwolfA5XFWKlmj+UGP1Aucw+lxqo4W6
C7xl46l0ov20ikeRSl7ZR3v+AThltDrn1UocaGfrGRBqEk6kvmo/7itEndT6btVxy9ddjTrHkoVV
OVN7yn5pzEsiHdapA04xAOwIXIGXAvCz+YwUxPXfLUCLeE0yHR0RLdDBBHNrwmsAo7rMaurkDN1o
F5ufw8XSsCnU/rF9jKIVGdG7W2HIJpiEFvpH+8yHTQSoOtZt+TDhiHAMC/fxKdZ0kiQIRDwjP2BZ
xwwYEFS4cToZQyTsIYOK0EkFIncuYmjzXojec/eVpy4Hr0xZW/gSjL4KPNTPPywEpg0KC+k46AYr
QqxAe43eHdzSDvv3IbzlhNltfvWCl1+Pw4IS1VsDYAkQmsre55lKpkqz1ZH05DQhX1LC4lLpfHK5
y/fyTN7NYnwY6M/IdjzXZZX+NSSGpCJAEh0+nA+rRXzVpREh5mJ5D5u7cXEG00XZBZdo2mHFI7Lz
smW69f+8ddSIC8UDx1Pw4MSP55nfzeOKNVUzKLOou+WJ3Mb0O0h5kIJhP4ZHSpKTfEvVmE0b3jBp
5xAB/yuL7YQivv7WwQ5ph4T7TT83uTedMcCuNj8ql3Uu1ASWbm07ocp5mvueIECLqdilsE0zHKHX
n76AgfR/xNAVJRIMHbzSG+o+TsF5oZnVcJw228k+oyWqkFz4xe+8uPBbQlNCpTS3e6Fc6ijHx9XA
kDE23E8UvbMLmd2NCJc8K8Fr3Iee/6kyWpm5+jSfM4uINxs7aDwc0OIrmG+OTgV4LwOxHPbmrxS7
/NwU0lYKJtFDBlg8ZpvRitLG3M3HvrLK8PWkcBAdq0srGpLNc4g/54CaszLXt5CxX35+h0KmtZFS
ujsO2WllYA+hzWtjJvOPQl99JAwhpgWbEp6YWPGwxw8yhz6jb5SpjsGWwyZCjr5Tw3yBJKrlBv+m
KTFzcKCVQrrypscpsU/8zRmKEetMpNVQhbKfQvpbNBNTkoF6fWKgUQGeoQf60j7QWZ94SAXhsuhl
PlqkYborA783uKlZr7Z91l8Vk0sijW7uTRSGoAlOWZDr6MO+hjOcN6Cw+bULYvRkNwsSNz2QXdvk
bhUSLk0q61gLQ3smL1Y4KVvdEEX2Cin0WVtRHaZHIN/aRaybueP6uBZCi8fhcuilOlMIeTWHBCK5
N5lcTyRuln/NZ8ydO8vPqCDBOWXG+oK5Aqr4/swIzidnoSwy/Go92EIr/csM6WAPp83WZEAarSjs
jmb5YYmLyKSkF3eXseSFkxgJdMbEOP8BkL5ObR/ThqdUfvV3OHRTfNeVW9DlaRpRRLOS3b/ix3+8
hYNhN9FYFobjflrMplgkVrGZ9wvb0xMbSvcSEu7EJGn4mHOTURDZepmN0RjqdkQZx2/T4Tt4sHgW
MQ0hgCA4Z2g/cKCw/jySsZ0op4eB3vT6G5LIciY9X+VE+YGqolfOEzvKcEmH8sK7QqhVJoHnRVlh
wvWF5v8DBRGLu2WsUe+O8tEJW1AwQEUxZhzp1LN3Ks/xaU+zwhhIVGqQwfzYW4T2h+Qjs+19e+vg
VpO5VKX6BOKu8cYXTFWbox9cfV4TyWPD9ShuuoJ2geZcXm2Zr0OiUVyKOLbA0XaT3ERYt5bcD49L
pYtGXixHVLUXXi/4c6lNmhQopxoeIqEyo7Xo7/izLf2IZK4ZxR+0b7VH7GvFHsVfMHZxU8B5vrC0
MMOb16VUVyICdI6OpmmdFCBJFwwnPqRJuk39QCA8DW9y6ynHp4Tz2LYXLh3BvzYju5ywPSYih3UB
mB6/Lw8XjqdPUkT5NgACNpjcOIVPP2mxDJU1mWu48hClMk3all7C71BmnQt4c70dEah8rrPzZt5R
ER6FsNkWbZUHZM95FDA0//SY/K7UiHJ/HyqiH5No4TBHuiMf/wkkuv1LZMHEA1uVkiR1kfi2PUyk
1efnd9clHfAOBhmzZ7TWVTSnnEMWxt8s8aY5bVy+AzcziWOkKEhDr9LJLDJ3Gr1/7zWcXe1OtRuV
ikilqnJw/OX4ocB/9Yx1eB8ahpA3Ckn50e5i9EagHm4URv+EwJQtMC3u8JZCmvedexCfmtiVAXjc
BNTfRWNXFNSZbWhywzTXmPZSQAe+bm64LYIwwx0XLiKdzfu9sichA2lWx+5Qp/Fv04s2STNuMmRe
3+8ztWbGrotHR8nCbmZpqCSHBaYdF4lFoa1lzEa6pe0Tlfgbe7U4b/gR8zCefN1nK4skMYy3WM6Y
YdQAOOeBFpPv5md6EhOWQ4u+oFqIW8lDIsum0q9ymmtUjgGR0WfE3n4FROj5VbTc+0r6wHe03m05
OPziXrpn26zrew4chkKAe9Pvu5wmu8NrNLaxLRASuQxNJf2/GwHg5YFmJxmw2JrCpQu8H+yeONi1
Lo7Qo68+MR7+R2VA91BdDn3wsYlWNCrJz7OZllIx643o8zYB+0bJowakzO4EeqX1c350zA8lTezD
wR7xMavAGY265YKjsbp9lGFd4kTLcC+2KFEzjyKVP4RmL8vrdWaCxk2rJimszxRxc0bEPA5AjpGR
J+ukqhve8tYpvI5Pm290tRYPf0hVqmBx9K1qOUnuQl2i6UoR82BSpXp2KBdw6nswyBcGuW093KDj
4Qj6uakUx2l8bwKHF+X4tA6M706vTLL7OrB1NQpmNkpB0SHRzo9Wgo7G5xU+ZDanKx0Pz4ZcGDqR
OWYeFSIXsT/2kU4BEszFe/08JZDgf+x1gZxEF8Kwej9YJbIMu366MGTP5yI53AjpCHhudHRrMhcl
Z0GWODhzG6iMkkXjp3xeLaV9jCB7/Rai/hPuLgpJFAkJIxTFnxOqHXrqwK5OMcIOBpG2Ngyq/e07
6ZzJ1zf5niHpufj+bvbKXbbsD6sZ3ikyzDyMnQEc1nmMeTZoZQZjTsVsNSPXnq5B2T3oZPv6n59J
3AGxc0GzRDDsCo+kR4O7Rr6eaCvFdwwQvfLjMzcGRb++1bi5ESLDdZ08GH9kU+frb74l2zac/L+y
rfX4CfvAWMpGCSZj1xlCKjsu13FOT/wQYk/ckwBZzhpTcLj/H+fTXuVGEj18AdHab+CyibI0tB9x
s7IJrY5EatxQ4mnpio8uH5B8dd3FqdrwZWnTgttZbWvwqEHRlpGO7Du9Wf388k4hhzGmekYFUHRk
6OXNTV1/IdKZ3MGHZ3y+ykY3RHgjyYGTfS0nDhN/ZngPv6CHynPuBn4161EXI1Thr+5ZmQI6D4Co
9YJahXz0gGBo0f2AJawR72loM5tuh+WMbscbJ6PW5VRHO4SPxVzfTDzFmwuWMlpiPEFAEUmrlURE
QZLVLst3V8zSzNsZZ9PtBPoMNc8WAZeuDnlm7mevFla22ryQPdAHiRZldsgx0IpCqn8aBvUYEBC/
FanHOfVRQpJIywnkBYLaukltWtyPnlIoq58qIhTUZSSkHtX2PyVPqmU4C2OfFw9xb7wLf9axbBiu
3Kj4vJTCid7iervA/wUG7F0mLjBfz3FG/JAllTJInC5zSWozmT5X0J11uFrvKWcJu1U5Cwk+JSx8
klFiP3CzY22chn9kNvMIj6bYL5xi96S/tpeqvMEvrhyrHVLA13OdIuU2StLRVM0/g4p9J+fAVJec
pe/LVX86fmdt0e291alNvv3rkgcctduD83t2MB/zQNHhp9oGdW62qRmfGxoaS6/CPlJvq5Ed31KB
g7vl5frO8pUIIZhtbNUijqcGh7eHQK5FOJxCGO8RYhmJaGcPAKBAu6SAj1DeiA+vqRnfufEKBi/7
tyfnCbMwd6ZD70fs8lE+ueAcd/aXp+uig+cOJ9TFvBd1loinVECL159vJehQtY5/grFwTs8bozUQ
Oze94Yb8r3Syd+CYBc+nkDf3okZxJqhPYsyc+J/OzqBDNCzCbanODP6vUL+TzlpM6tpJdc9uBDaC
oelVeamvOVHdcGyqTw8nGIf4L3lNy3t96oYaPcfiW9dbVPSxcRP6HYUPA1/4U7+vP2tssuoAa5kz
TYgadtA7w7lkTm4v2fWEhrrw5c7wkQ2yl4VqpB+3FZmr9XHQeb0rsZYzDfkQIOQipyCwznBM9Iyy
2BjlLLF5pXPXnT87hPzqKQmWUkhlieJWhW/DqDq4F9SoDrNBIKyDC/6MxxzO1RTAJ7E8gZqYG6Hp
LSr5cowHu42NiEUWVp/gTvM596PUqTBKsuxHdOSHaI2bxYZqP4MRFHoRj4KVzZUDIDVHlDs9Uwo9
u5XEjs3hRyocZ8/nnPB0+ED+NDbpPbZbxGhg2QMDQ7D0jaVtNIQpeOSsvkfUwKw7bhrGWlgLNQDj
lMR0zJb9s205FwiPD4VcPF6dbRk4517ScMj2h0Bq5tEPUFZFzWtdNFqvDudDxW9ykHNQMl2yMj7f
REIRmlJjItbFQJLkIJlBXrTxXEqKhv9vm+ziSuvTWJbyfIi6XM6fcBsujgEAusii6sS6ZRDe8RTg
cmC4NSAqThuG1MQOHyL7SFnF04MpuC0sONop6uKa7luhkZ6JUUJi6ARVwXoHcntsSEIwF4GDMRNf
mvI8Nfwsw6eSAESdLmVTNPhrHzRCf3BbQWTZFB8H29cBE/Ka+N1pHqn7k4vE5jpxhf0TLnnWCKho
jRdQ0+kWQuELInSVrnN2TAR6zAYGazf0BOw7MGrYflXoMQV2bJIzZuT2c6Hj5rmAAd5lI6vw8PI/
IK3368VD4crzpXhGayOtEU2lLDRjCy3WhGAILGgesq81tosahvABrSG8nIwFNavNXvrh+DyD+0xB
Ww1lrzgZCbCKiPtl2d5xWCtlwg9K0TtTnz3v/mM4RTV3qFwUxoAR6tjBkBs8XCnQCUei7mMghDIn
Jo8HqPy+v0XGIJvg5Bse3kdovgEfSrTug4tr8h8xlkyxDw79qdJjaTmmiBYxvqqWTPgT1m0bXKF5
aCP+6BnXfH0Mr1duJkUfoIwf1YWeZyc8I7x1oCdVym/4CCZP44hX/LiWur0DYg06XqMaH3IHBiuN
YZDzW/RPX2q5ov3AWW/eWJTodsMubh4Z8HJDVRbXwGll9Ia1Jdxbra6KAMuGvN6X80gig4ObcYBF
tNyPUCzBtYcQJ6UdfXIU2BMipk8HejQVzoxaFoj1q8X3xjVSsnyLP603DlOjTCNjVuUYr1uKSS7U
CM2HOxDZvT1chPl+6qt7iJVuey6IrCnTRgmnJ5rh0XMbDJ6c5OeX1PgHylakZfXi+6jUPui+F+24
kUyCgJq/l+mhS0qEaW6GrnkbH4omvdo//wX6BqLXaL03XrnZoDo+vYzsEasbCpbqwtACnwgvzdU4
tmu1Ru4IYlQfy9KkbvostSWP/VpMUUPnvzpFeLAynGyKSbLwtk1xeOuumHEgWDVd20d/sx+CYFDY
MWjBWAYD2cFsziFqQHK+UIGZf6hk3JSqVtmbHdkqBZqqtyLvBQ9WH9NwrzKlxtY9KCZhbx6kvZxQ
YOtdBW/vaYsv/PbczKwcKYQejW1HrpzFc1Fz/gBDkT5jXmpDXQr1aBgw8qvJ+tzNLXvYaUVGijkh
6oadiG0ExCbkuv5px1/9aFImczeZrLM7CkEoLuQuZq770KiOCNesMCB0AseVw1HqXEz8ynmT744i
TwpksyceVGv4of6rmZLGQrHbp2/9IVTpjAJjUOlSo1DfSOORp7ykh/xAs68dvc1VqIz9iC30gGVL
kAz6C06C/ZvbSB9DvrPT/yNJ7MlRxY+HXkCZaQGqcO4RqqyeO6BBSi354wdbtfQUuhdy43pxfwwB
wdWl+5DnQVCViqkcLu5UhVGEMjBpTQbE4RMch71LwxXNisS8PG+3oGTayb0E60GYxG+AoYeqS0jQ
gTDaQ8WF4aii+CwyouPtwaCgRP8klpO67hI/oakDtAVMaZbfz2iAT+woHtGwaey3dVZcPsl3yezq
Qucud8bDmIeC3Ufi7j74KMn+6aOtezRKXZUPeuSpD66WkYQZAsLijokUYidtCPydXtXEhgK0EXrQ
ClZhgqZlcsK2K6DJbfjbr5lLsmPGSM9Lq3854OH4sPmFioCYuHhNuR2Wd7hJcOWMpXAUGvMWON0s
yCsU9XCkjJqi/53ZjlNIe1rWIv63HYZHruQ5TPx8KRzIMFoLLGkMDsMj/NddQKYDai5bfidC0N6S
dkhZOQyw3rnmDEKbBOdkgQya1Ec29C6KRV6x4nsvZmZHDMdns71njLbd6jOK1nuXdTz9cN8IQ2H7
/45EDL6aQwE9Mzz5z9lUvbp/Q7Me+y8lcTbrJengftq7NJlIdOMVvUO2CIzSBxzou9WzV16EViu3
PSyFlshqgRfQNYqzW7CZyyf6oCnotAzhqOSKCk2dXdFgaGfGfc/WjpyH2Eey0Zhn40ZXEDVp9DKe
T/GTBnBMrjHnE05f3EqeSiRYrKHAx4yQChWklYFeN13mo+tPuFPHAPg5W3LUVv+tN99to0bOynyW
DA61eJ5vnZeRXSbocW3bVFIWy67cDCOrnedNvsgY3J/YFblDFnxxy19phsXt/l/g4wrBdfRLwfrL
JKoUEvNLmqWHVcvZ3cNg4wjcoIR6WyBfHnx1GBSKfNbXpf9rASBzXIxIKbuy6sMlyn0LT3EvWUS0
cLcG+uLu6c48fvAdBu2D31bFfGU04/UT9tAp4453mVM0aZzLZ9lTOLnQT6JRLFA7zH3OBm056BT+
YfcWWGG992CW12WFBvmruzHEo6DJGZ7TrmaUKobAtFGohrIJRZYq8WsMTXUEC5sGbozP9TorVN4I
TpXmyoZePmc9d2xFfqa7tYzh9cNIIHYXUoRRSSti67WCiTJ1EBUmo6vqf8F40NeBbhExJCV0mtUg
L1GXDw3xGahgZK0g8VOaZFxlVb7J+OInLspNgETeU4HhDxOpnX4HfU67VSSLqDKlgFbLMkQD+/U7
DyVrawJ3gsVKck3Kfy/ncRifVnlqvv3WZGnPsN1YhY2W0kJuKhxKoEikPngLrkd/z2ZgIpxYKLHP
UB8ll+q5bMweFsPDYCCgFY/+ZpSbvzoO1AVRyxkFf5ehdNQb3CGpNNlMyS1yElqNQgTwT7jfbqiC
4qWIxuL/WxiBOqkgyA3sDs5hh814xZIYeJeKnM+hoDcC9Rg9zHfzH5FP/xOPHUqHWmc1r0Hna7aq
YEa7VqIVoDghY52B3N3fBSHS9BA83mqusHQBjnWOra7xfWvvrDEWqASSON5QzMpArcaL3Gpz/N5k
gygGZyP3G+o147L/onfLWZyK7ySics6/yrL8IqcH56gusB/m7ey1h/tlmLM9hYnpPvbOcXCbcfl8
yey4X5SHFboVdIgRZh7yfxK+mOM8Z68VPwKGZc0KpLseHcRgWSCo/IG7LqMNXBmI3MsK8cNaoHaN
fKkeLobxcXKEk5O53YruRiEkHC9FppkuktuZp8/j7NCoGsDipW1LhJwuWvM+IebkXzxKEZe+PAQa
pifT5QzWluFt9E06I9EPX+UJ5FNkAvyhaKktHCeoM4T4bsYDLt+1rIplXDmczQGSYWLSeIRMbAQC
gDTJhrQWmAAF5RbgsEhkamNdEJoQy2vLBBwijf/eeq7xvvDs765pC1xEnVd3NtSymOmjIUwSHYOE
prAYf0dhzNDSl0bhmVWcN3b73AqzjVu4yEaChNFiE6qCZoT64KhGDrfpl7VbgOYj2gWILVkfZOh1
W4+Jvk19l0G4Aiul9069yLSyzD+HV4kkijdlxroDRhwymAG9Onkwp6Nv+gIu37TN/qE+K3IOxnv0
yr12njS8QwmW4+XupKQEzr7K1tXdxFuEft2q6wxu+wN9GezeB3PZGmwN/sOmSRLot8V5w5AJh1LC
03iwU7fsKMXRJTwzA2aJzJj9Gfom1ZRGOpFdGl+WDYnVKmOdpkzd5xQtn2dyrhlFVNdnlWbG03cW
F6ebno1/wWZXnRofcpdNYGMPCd0xYYbs7QfLphndcRnClT8hGUB+lGHI0Udup/LDK224DN5OgZEd
7uc8aTXCLNc0KL48Wn76anureKnigxTgg+LOkRe4hmWwcqcDGHAK4gnJX6UALLj+KhFn+b89Y4FX
TAdsR7v8qFrdhx2pFEurbjr9i+Q6tyrcs0xV76z/RmjLn/zU6bMGIB7n5eKbpPlWuiMfjAEGWIpu
ghEFGcD9VQd7/QoMSBZyjS8E5zCbvm4eBK769Fdbc6ZJhwM4CxkVKmUwkF55Gy7TEQ+bfHy/rvVk
uCCrgYN/VGRcJ5H9hbZkHpduaAw5GYc6vFXEFd/A/UPWy86F+FzOGWI3WVVuA+Ymu/4w3feSRX4/
4mYzgjPTkeKlJIHozfjqcPQqF4nFTSo/HDdEWMBhCThJhgveoKQakv0Jwc8Or+5yFQaJnwm2eZWw
OVRpXMO7+38d7PA/lSP3TI5EeNXl5bLXyPWYpsftV3I=
`pragma protect end_protected
