// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W/g46+5OqzLI8lmbdzTg9cbtiRMFf851hVFKLK/qOm3jWD8FqVoifbAPYPo1Txhu
0pjZR7+9rXC15058nMxjJCKONUOHJst6Qbk3Ce6cY37+XE4imeq0vgbvQjDZI9kL
SkhXo8KAHje79yhwJHGIRV8TZ4fItJkDz0ESM+4tXa8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
ZPxh6Ut4YBFKZ7tNpG3RzgWakYRdKUMXisbqIrbE/3ldSgnHWkxpuByP/g4Hg0Zg
TFAPFCSLNWXvsSiMm67+pzmR4CUeeaNAtvpeTJpQmM5rs5599urtqSgwOo6PjYOl
hEE2gMRxp29XRcjQ0F6A8IlEPL7iXc4apajaPKkYRA125xSd5L1SHRbZkbE0A65l
SW1rlKPrNsdVjHTCaNUrER8UwuAjW4O2GFil6TmZ6S62kOil/thr7JcPzl4SjFWN
DkqXeOCDsMXp7XJRrJ1iH+udOF22hTenfnZfwX/BwYdE9aCwKJF+VFJOkuSii+v4
zDKJyar2IzC9MrOwAVp9o8axH3NStLAdtizs36V2Y94lU3VtSWMxfjZSRISuTwSD
Bvq9oanVF63ZyrhHW0jXNKumJ48iupLVs+2+vguDZJ+LJqX+tvXzquPsYXtqnGRz
+AM8O8unGrHZDeog5xuWXRzrReXmCj2vpUl68sbX/ioqJxrzs1HV//cu81b302rL
LDKYQGIKt/AIKzZ9w5EyuaNA4vmg+10gkRsliPVq2nPfLivYaC4Rw/OxCN7OsWO3
Id9XevK6OO7rmKlh+glSHC0GLnLYg176DMFUa/ERpi0Tm1gk1j2OHteAPDb1uNGA
Lcwu02bQZwy3EwC8rLpTfjdtHYYqkag4xHrGt72drjfNm8sDDbGnmL/3vdgFyroH
bZ1RETxtUAs7fGYXjO01ZWigB1jm6qa0qMoryNaQ8rSeChaydMwnHeYkbid37EzU
zK8JD6GJunFuLHGQd2xiPCOyW0boNXJ7/GVHsyVKiLN8rKOXlPxx0BrK2tuwhff9
Hav9WhFAAM8+6ffJEF9GIX7wo5BgXzJRd6VvQA7CPd3Y8b/ydJ//rfYJhPQQIcR5
jHLDhRRuYiT4yCqPUO81RrsLZFfUTzehd31iZUZdQH9Wi1AF+gU30CqZnfhiwDq1
D0E6POBiSd982IPOqRKYEZZIfz2GHEu0fn3+cHfqEkkUKNDoh3pxFi/KEYwgYsNi
/mvfwCK1dJ1WdFiZl08NxiyKO9ad66nPamKPxdKPqxE1jdy2iMe6xOWen/gfylOt
T/a6godGjL2agCQ8F7rJCJHw1PttQENCBLZWT3fLGQnxcUMQTHb1CIWfuEUHdzMI
67RY1uzV75OOdPXcTfTIVvYcnjEEvOHPMnA3Qbc0Oq8qZK+2Qoqs3gry8w8Tl/7p
UXcGgvSkp7gs0I1ggJj9jIsBEpTyevbWiVw5pHD/YJwDSjZq6AMIBqkW/ATnGIZU
dJJRKQ5IgVVvy6P8kHyzIdm5sYmK0heYl1f8Cp/+B+C+2p3igj8eSmQL/OJ2NdB0
R2d0VZJoxg0JkWpffcolhg5gyUNYMwdu3aUvcNclKe8hB7BCVuddPa1ieM0mZce8
uceoUUW/14mi743Z3t6Qs2l5qaZs3IDZCMXFSGLY4QhFU3KqmCwChp/ZjW2FhA4p
3YMqE5KKKrxCdK82vkOiItFA2NmPbXB+iyf4zkknBn5imCpr9HrnrS6SufIWyLf9
0NteCs0Fbir+3WWSOL1zfDGHQQq7O2YX4FLH6BzkQW2wIvhcbUGC01jaTIs69Lrt
ckA6VQaQO5eYbOEolG1hQrib6YLBl5oeez6bEwnnYcvaCMHlGQpmIuqQuAWwo7Kb
Nelmi8iL3d8Y87EpWiomDBj3i/TFw9x4hUmgPphpspkW00l2Ca6MNn9CxFef8y+C
pify5pnOrZcnNvzZv5wwU1paYAUX/uTjWE9O4sgmBEkXPy+XfX5OoydfCiTAe4rA
tosrp+m8MnZHzzTkil0aLMRFbItRFhMtBBj4H8Ik9zG9nVd3mkZezlk/btgPPK7n
DQz5lYnumEJpqjpvGcVAeXHUgBrC7WLD3IJ7SwR2OchBi9d/CAaK4yvtdaM3VHTf
TCRyvLBSTTYFpNpx0Hu5VOrGzPXfgo7iY509bUgM5wAYdQ0+O/IJ7U0X13w+YS5H
c0c6YRoHBOOwP07Lrg8ZXRHD6dHvOoCo1mT23Jjd26R31p/ChdAp8AfOOS6EIHHf
gu8kJGH3y6W+OxlKdaSqgN4jfLmivjOqr6lzc97ehZlnZ8fDqEFSSc75wS2kUiOy
0yu3VGeZS19cdmFI26qFM+GBw4PpPDvxVYiRimNpmKWVEjo8gJuyg6k0UZNJgkF0
p80+dE8tn+qRpATkRj0f47JCb5KNhaB6zv8HC9TAAxz+5o7WHHZJsvbAe1zBzITk
beFLT9SA94M/gKpDBJHFqw80jfg9qhQRFT9LRE9oEuXVc7zBBPoM7G1iLYdWMi0e
w4xWW7jkXZXOMGluFTPbEB5fZ3sandFXWMJRofgGEdj0ytCSbIvuTp5Urd9+PPA3
AEYVTjX6ymUfOEs3VnScI/4p3zWWqwJO145d9n2/eqO9DFlT6ldkBDJWlWgPu07j
Pm1YCvbBLnv0haraEVcZxs9UNTgyhI/OzN4ntgCY3u6NUj9n2Jwy3u8Uv1FNpDL2
VvqIqXxXmw12wRdTJw0u8KTZbBiJvcGLJw9Ggt0/8eq6PiRQaOmwA77lUhYf7xN/
rcDGXcYHyh936Qt/leVwd/G6oEcOOq1q12s2u6bnnhu4u8mzjUi7RM8mtshlYMij
vhOKV7Qa4HT8UC3YnzGnt+5EG2DqOGj9KI7JlC73djIae0T+MqQ0PytnGdRdDGlc
0ba9lvwPfaoN26Uf3FkRPrHcfW8EkEadZgWk2fhadbYSOhjrAAGX6pmS43kKw/xT
9XEMielWkjMKTyZYdOa6RjYHtMYfZ3xUVlRE48Qty7opUtw3ypND88/0Tkoz92+d
JSeuoVr4GhIhKjRSHSbfz6fg36/lqvWX+KCk59LPezNEqxRSdCmK7yhGFyYbWTUO
QOp5n4RxGsrFhO9aWgFCuPCISpcLZ9z5xuMQsMOpQTxeBhW4Knre4B4LpK1Esx/E
KmAxkkeSgdczdIxr74DY5448FFKI3zfp5dj3IJvEP7qQzIG4H/sWKX3IL7/pHCAc
+RRonueBown3Q8MxscdSwyUTIW1mAj+Vtp7MJVlQAEOs4ExZ9WK4o/yO9Odr0WRz
ezVJZuZBtGxSBL6FBauTUn13Ujm0+kTq5XeEoK87mkfsQ/LJ1SCCkcTtI9RxZTnN
Hce5UGiZ83KGO6ZvfIEZ5yhnAULwAWX9GHZ/6kiTfg7rAY18JEL0W+Y3vPCBfvSL
/KEsOF2uNupPaLtNk3uAqcCt/ZLCIInWKmONKDfy3kCdDNwNQa1RODmdN0v8prRy
IERCgNMVddIimBSiBF9h24oGziQKubGtnfiWl2mOt8/sNfxbPQRqLSayupeGbEtT
EdaBDSbnzobVWiLMz/qGXhLW43Gey+7BagbGdx7aoVfqbz3tu6dKV3M4kWzhZ+iB
bOrsNFV6J7YyV+O1xFR/3047aDuZRVf52sv+CsUkbY8V7hL0iy/nFOT6xYHsxaOu
YJH52hVPHPjpRimHwUw1Cjx2J1WW3kcbx3TW+t/qv9ILR+lpalLLgnU5VUQlD/4p
pNAG7C3L7/XpK43FDtIrzUFL8cNpExdlDY/sNfovW3P2BvdBojbVvcPe0gdyHWjm
LI61tKxMgYSqZCayFOxj0Qb+rRQnFnU9EUZpZYWnYowH3htqvYZJ9C09ZpPAbEFz
0BNeTKtBgX9Pqsidh1vNv7QpjiN2A2MvcC7BFJ7J+1xzL72c4XcbQupe3HI8t3JD
X6v9/0jn5cYL8BqZ+zKIh2CcRFKzlkcL92Khjwv5sXyWXs3w2zwxtTwq4e4SrhBP
sJK4w9lPcyGvVjqkSSdjUNKaST9aqxZ/6Eq0sfRFtP5dkraPmO2P3SjxUst84+jB
Ulf5Zsna6gZLBOV1Buqnx8yYRCVcdeRTq5nQeZpqU11zEs2AJdEHXjHp42gOGK3o
Weh9dYPrSj7agvOjn52tNOY1iB06+hN7OjdaJ4M5XTWW8rRJTnysHF1DkcD9Dt6d
MVyACbl7YkSXnyPzHUY1Kmgaz0V2SCjUuc6Z8iB8/7tEUBjSkiPMBMYY9gOPHb9o
/5eGxxGP5UNkKTXcbD2Q2keerNjPIEK+n0RXgpTxpn1P14ILG840M16DSqPbpzxn
l02Vu4YgY+RpH5VJw0fGl/vkwXuO3gRnSbbb4QTJsUpUmNvvgZVY1DIitrBShZww
uMwWEEN7SHWG/fNo1ffHply7jbjpc9whCpDxRQCDqZS9E+47QpO5Vfa5IFqxlZLs
GqJ4f96k/GEEx+6auC1e923ekZXEIzBy4W8n4qBloaA+wtGoDKDLeLP+GoCJuQQj
p3RoYbqlZ37ZmNUu3wD7QG6bDvGEk9qg7doGemxO9R37C54YvYgguxVbo9MVY9jW
5tcH5hx+xbYDUACZ5D9xNUvOv3fXjsDBS+XcjRioqPZTS1PrkD5mcu3ledywU7/r
MDrH9A9BpIlTlrNU88PlLv5FAN50dKdeOoU9y3xpNUeFIE0wAYz2q3pqDGSa6leo
lexTXIPVOtswtvOKsZJ1s+w3qwrR3L6TUmOfJSNHNTaoLTXWEv3T0QjB79+VXbOk
2vOrBKxO3dlgJlFD3on4BP1HMIKcRvidBxwA9+hltegYNXivCIg5HyXFrie5kkov
/1v7JaShGdWf6C69ze7JDg78Nzv7tDCeQ9wnyKDQVEH/2fjefFGdoXrx/De2uyiu
MYANGM1NG51Hi1JgzOrTBduG+TUIK8bBKGSRSexOPSXeuRrB/MvJ4DpvT31ZsAlL
sL/NiDOmIntvCw737GIukiftX5qtOru+nAj+ReUKiQ+MiMZKZeiypS+F/rBhNwkt
1Td5cO3b+bkEynExchq35+H9HxJrYTYIc57V9bn3eD9RKt0+HnYRrDCwh1NckBbH
6v2oGCtTX7/+A0ousg1TMOsJvButRf844oBPl7ke4c3fO1iiyfzICqSPNhwyRbzm
mfLM/VfSuORdHQpEerQDapsypU3sdeFfEk+AsYhm/HUVHRr2U7EVOaBlHZVMK9QK
XXOIiEdMa4FqtQ9y8V++VCFSOlSYseb5RpFHrVU+ceUp1ezDBOHxXUkyK/zlrTXx
sX8v3uP5Y0YxJP/UcXEABDMQIvjZCLfvS1VuoZybDFesA2zQegZ7ETZjo36rUM4S
8q31kruF69BGlvpDBZ3e8u2aPgy1IEbGyTw0vYWuUJJ02ku9Ir5xpDTWV+YJsXwl
bg9EBufT/obE43rf0dNVKd5iS0nNCM5nPAIVlHxLGv9YPW7KQE/NAOyzvQk/j1Vu
jU9nkxGtI3gQi+A+QHWbvZJsJTjelFX+m9qjSuLDiNkibGn4PL1K5xb8BGUWvc70
wawwNFjtakoF5s0ydiu96xKHLmf9yeQPJiaJfBTDWvXhE0SboN1J+iiEyqZnaJfX
tiLSLlYHspV0XecGn3TG4dXeeRth3u3rR8pa9xTxwws2gyMH1io/w/IIbRHjMF7Q
d61b6lUrpb4LnS39+Ih6JmmbgzUwopkX5JbjSGgWQxb1LuLOWeTljhIIIaom4YwE
73AsIszNSNji3q3DhWzTzlqvZbIL6cxC8MW8X46roDfLr6csgQbk25b126Djcywa
944G7+OePpVlfoQ5OKNPEeYJaj7njuxMS7d5Lj6DNab6KE/N/qFfx5GXcUjQ5qss
WdB7XlPIBlTK8OVTeHFwKFtuMGgJjnz0JQFl8F6Kz+Aiw0t7vZJLhUKheq4KGXAu
ETZDwrDfb+CmAqwbV/yv2kGbirJYsbh94Qo8VGKHoGo9pcHyp97dymiMVn46gpMa
qjgTUf6iAzhBIx5m3rMbZkpwbyBeiKnbO0ZlRLE12HlQ7QI2qVKY+n5vMxhD+BkR
sV4wef/1RwFijRpg6gVM2TH8zd/axpYBlKuB/6SXlDYWX2DFxQHZY4/digKPb+O1
PbGr2Ltk3JZq2hJfmVq2WXdN8OhVpilxdmBTq1i13Mzlv/IXRzw9iK5/j9VYtGlh
Ei1CABCMVRJCHocppUB3rsGidZWjW5DYo4qQMazjd5Ugo1zrzfBeK/rSxBeS9WyJ
DM+0x90g4rHhhGCaakzLg9AgESqIekdaUHQHGk/CHunDfDjvu8Mlh+f3oL5466sY
UKzTkLhNG0YSWbXuwMeRgWulKp683CIBnCs764l22XaI10aH8IjuKxS5sxcsQskC
ZjTfB2FF0frgcZRPGUknbMG2JalBdbRDZ/bWy8aN9aEuZijWeHiwEOdp9VwIl1lV
AxwCFI6VRRUZb9gGCJhWxsuSfsR08K3MkOIBeFoaQ1fKpgfURreBl9SRVDmsRuwa
0VPsnJP/ZLqlPGbV4zFlP0khUjvKthrDhWomVqYxZjDAjCxZpgiKA8H/pisxDUKn
vy3N7Mkg43BWQHu9dVMpdOWijMqatZGqrQjTlqkSRXSunKZu1BkFocAnTeVMymbO
O78OUDCU2LucDbYg+36gN2t83FDKrrPGpv4Idjiqt9pSbAehyd7OJYBEpmRwGlwo
c7n8/Jf+52PUWYv9JJS46kwJxQvUXv3X6DAm7FM1NmXCP6Ro+KPiJMpFKM0+4XY+
RePQ/KZTdBJTPPBh5jw4Shc0kB/cfgIUHvyBQxqPl0q/2FTcHTBQuTEWNEQs4x//
h7eQHGP0o4nLZB0jNcSqIB1/NDg6UD0iWJrGCaiFZWAYQ0rkZYXR6Zn6W0KkZRIp
7FJ/tvZQtimnj0WdqBqzKthNV9Dah8eBV4RlO09XjjvnC0umZVxY2nJsnAd91nd8
bMwqiywc4TAfnw4H/7bgVzHawaFipKZYVG7K84DFVHGpeK5tKqlMsvlOzIlDUdTj
2FOtD1WMzYRdfAPnrpdZsp9Uli3ael0cPwx0il1W3990xIKsBo6r9szS96GKi1iJ
tsvywiMvw9RT3H4R1F0tsbrUcFqEW0b4h8omCf0NIrAB6euo9cKpOTM/5ELfyq7b
lWShFOlkC/zLCGEWyz5X4gdtmQe43b7f1kVYSpiInlj8X1PZIpO8UHxWEsL7d+VN
17KSDXBP92qaMHJ+yd9zlvo9kM4BDL/EH0bwEMVkYK7mIw7RXzBTlzVYElt6G9Gl
Z3tJhVEgLqLNnxk2hvxKdHfpN00CNFU6Ep6PdzIHS4/cWHYfgkBxFKCegVn/iHYP
64n92eVv9w9Nqg8N4DgzwIsE+A5h8t6Q1zMHTFMQcExXwwVxdBXbyfeiCeYfj2Zf
GYii9TogKlX52fiDOXpXdIC4/NPQrQDhakZF1SSB15UrWnVns30XPKlKFdYVSf/3
OdYcoyeUIQxvWIYRs/7Gzt9IzKkcIukzAijKCsBo+1k/kNaRyd2lAbSdrzGEcFnN
6IhNgjfDhdkmRYNdszW4uZaPaps0cCqEfhNSOVlnZOeHgPgu9bpXtCkLLLZeC7SM
RwdKpz7jPXV1asFQodNl/Y+hwQPalLshXMIH+aMbcduZsVFcI0CvDxLaDS8HZFCA
zmr334yOZUmC8HWmrkoVLTcfII7Nu/ZUFVSbVaLxTotbRSIFRwMtqoNfukXZXs8t
a8U9rTUsmIryfbpX516ZJMDHbE1uJRErAPDRSnnkxUR6hYC/5XvscQllc5sF9AaR
h8XV5444IRdU6Ca54FRw+FBFdAMYvSFeYR79Mrlbqtix+rRKrGE0YmEVxWzh+0QU
/IDHqu8Atd8vP4oXFQKBR15pMqXSDVgkAZ0i+skB+YSa1u4gXv8YCFykU8Oz2/6h
306qn9dQvGy2nP/LT4NldObdlL2rjEuCQFt3knkNuGkHLbjNJbDwfvKo0GPbE/Ne
JGU788vQBTiwk5IJdgr0DqS7tIKaeBYUaKKDqXqf3W4QA3rXSBz8kvyCVGe6VX+K
0Pd4TOxFN231C332KcTT/MAvctdCozTgUBIgxj08GLu5qcpHC5aNDOgdrtxftIJg
VduVO8QDUO8Zeb8ELGZtjYqKBmyFQ0KKhOxK+lPzeOnFv523TIAjAvHP6oxeTQg5
qkVD7t8uSHAhHdx3mtuUPxU92bSoRBU6Gt3jts32pmu4S7cmj1lFsHhzP8QyOQFP
5+CLbsqc86YeGczAUB5WZ1WLAEUmIy7/HXhn3c099sZlWqWxSgdwN7lgGgWeTlr7
oZmjdvKHl9Xfm3vVMmLfDpDBJppp57eYIxWMoiBKQ+WwM7+E0cUZkkM4/2EuuoL6
4VqXUN2v1LHl6GonmifzwAKf6Jwuwc2shnGzvK1k0Ywfi4CeZB+jU7sMWKxXEd5H
iTKgY3P2apoPUN63eMZO5HlUVnjBmekyzBmiRmF9r/VmmzqO/j0waZvpWUi61X/h
kuuZywDne14esgMi8jpGfVp9AdmxlWy91jjInZDBxVRnB+lgI+gA7GyH01Ro2+fN
vDkahqsQKYd80h0Yd84NJgAq1S7A7frKHxB1G8Evh2kDqEKZIvrpWof4IP33qD+y
u+stZxHXJlOjIAd3VlCGfRKwc3g0jooMUT0p190s7NKCP2bE23Fgh15yC7H3ANqJ
f504c2gFqU5Ic/S35ewwtbOdwIQg9doTlnXqPnD2VfpH25bd3vyDpRwgxIIdKRpZ
fE72TtT3q2Le1dWqAuyriNJhaZ/1YrVjmAJyTs5/4lV9xpfMw2OFzLO9YPQeuZo3
cDFNmmLkiwrXPaSOt/iRlpxTemKFl1S2ipvQCiKmGGNBij4BaRCPwDkYrbsp1jyy
VGLTEQ4LqpMsN9bxkuXGqkr4akzgAxqK2jeTbEamcnzHIQfzanYEy7WLF2ohMOCr
BrtacZ1niC7CqlVNt/ME6g1X7redHxjFWYoSxF6zYWgqN5OvDFvB36/5YbkCHcke
43oc3DADX3jBxHtWatU3TmNmsY5YrUv0g8G2P+vo0Bn8ndBPpYw8OgSmdF3EHk+I
oMpaPwqpBgiW8byWvgmQ1aPewgA02YSUd+6Ic+OT3esqZWUtuyF4nqAuHifMCB1B
73SBjl25WrODqEeQ+dj4gXEK9RQeSNAn39Sq0IxKL8IFmSjJXQTljsTCtjXZYzGX
BzYiPX+bXvyh77vbIrTSG2altjP+VwG0JoX4SwS86DoSaRjc/fGMGT3AYsvX5YQA
LA7Um3eIUldRtutnyFlEkEeEeeXOn9GFY8a91fzBUlmL7V2caOjKEHs+j5flYlZU
Tqt9gq8/SVmvMTBaRpRn+U408sWmyL4Axj5gqeOTeSbeizgGDdby6RFBIHhRbHsB
3UW5kUyosEL0DuO1Ybew5cpRaShv10qT8YxH/MQa9rN3l1TksghAHP3L2KdbpNe0
ogbUvpY+VZuAUO+hSBjJYu4PEW+qS/IvwopSQzlFgOBE7NrjZmXh9ZkGRQEynDOn
Ij/gXL3mvfVuhqZ7vKyWjtY9E7JZhycyPmOIJjYT52mXCnDe3cQ36d5KpTtDxxVG
U14nsDMoks3KzHrfK7rbbyftFli4bbIP3J5op5R3t6qj0oSKp2J6fG4u9fUmnUed
/Ocjs0sPG0FhOiDyMs2RfVknM7esfgkpKrhUrGw4AT39fbutiSg7zAs0MXWe5hBW
vJLWaA3r9UdzfLpWCJGQRRts+zdiZyBadzNGlGwPMHQLwr1qTKLBJgEh8MDa1oyF
3EfFshZHjydVJCIYgLPoVgNuCZn6x5SaSKBm/AUfmd7j99o3kcw9Mgg9BcUDGxmI
eUVpLu/vJsDzj6BfnOv4Hl3m4e96VC2MMjn0rEDSXIlVCcf6x2Ji+C0hG3/GGe+Q
RVN+V4vgG4mrUibyZ0fz0hPTBeiotoXzQtczfzmeCZ7SoDuxDbttGuf7yh8qLW5f
QIYeX3AUALQC9u2E/JyUAzDDhG2GlRpqhwV/JAjB1rRMuJ7k0nTtQOGrgnuGG9nc
DXCSpsoshWXlpV51B147LUI9N0w9s41G0xvE7sqBbdcyyHpr4MdwTLJnVE8Y8S26
9SHKAQ/mv0/xVKc97ooUrM1z3NI4eo1KuILIZWwzpRRqSW9RCf08ZdZWzVoHPD4S
xn6ZjUAyWkcmBkKmX3O8N7LpYddzsteSe7b4vMA8a9t2URvCUTDhIrR1J+5LrEQh
B3Xdka3tS7OZQg+A/ygZGyaoqOjGXX49MWYZmMdXxhbJfPsg4rUT2qHDbAhm1Zb+
Jb4BoRPo9XqxBkIY9bN8AxM8dRIAJ8cip8otJCJErcRG/TC+OOC3dC1e75og8Xdg
j7QVtGR13UVU/yKcIi5EBblhaOs3AV0i8rYiltjPUfldVtnR0tSkYnybu34YGVqL
SGhXUEJnlssPpUJzFG+/YwKm0XbpjA+zSxLXtOTakn9u0dxBBzLu9uo8iiPItJb3
X1Z5jBjKOBjY8zUA+986ka2MMCyFqodpBvBBiiFUucMIcXKM6nmfxLIwpwIjGtPS
0ousQB6D3UADgf4uIp2D8a19z77OV+os+yDC3Xh9iEF/5AL0VH2qZK/kM3ki4VKD
vj8l98KnLhLjv3hDB7cFAmUCDmCVWPkNL7Q5FUwjYiRQGXDn0KYtQ195N5WSgFUe
n/JFtzfq+4Akg/mwa5cGiea+ZJZ9kzdq4aGZTsEVXPel1ztzzuQK6SqSbLH7M/c9
r2cafVZTu9zfzHlfZw/DFsxj9ZnaOZFlV4yXM6/ZgTAfPUeNyghpn8QvMSEDDMP2
14GZmx7MOxp/tcvhGFgj/jpgXAhrCCCastGBB1RkW4hTpqvjKiG1I/kJV2h5N0+G
4/I7y8FbsWXtO4l57d3KMqwrESmj0dEYh1hdKjAgyuMO0wfsWp4c9jtaKKhSyuNr
uGflDSP0pRTj7zURKH6ekRnzAmUxNzGvK+w2Auv8f9mixvRqBPShiWg66UKGQmPO
c/S+IKp8T7ZT51+MT9NS62CCHfFYpzfPO6lJ4M3d7jkq19pSZ8iJXltdSGVaLmMW
767sEQ6nh1p7hM3lHpVzzMmxTLnUxc1Emguo7v2p6MCNxwYU8JsdJCSE4gWNt2Kj
fUH15kE7wduhokv9dBEkzLVui6qhFrT+Cnc60IOpz7463CFdNC5l5FDv21cyh3KR
WUyCYKjD1es1OEwGcz0UrW1rNowx373RhgSzR4slISc60NCCbL6MpPJxdH0d6Lam
AB56EoXD8m8SyH1j7FiD3p2ibYlYWHy4lnPY6QECCdiQ+TTI0AgVqyuuVO9E3snN
PPBrNE1n5Ek3abEI/VQxHfg4dmkMHH9hTWKcPM2lcJLLnFwZN3opXkdUDwJEOtL9
aU0MM6oIDEFA0NDMyTZjTwz6QFX/qYSsz2sm6RUM9MP9RxSG1sUeYzs8lt2B7wMk
nZCgFiDHB5+iBbx73Qg9gLO9NyLu/AbT6FFmUSQOJwqGznUvTzzceSBYmHxgCEOJ
KjbmEEBPgLANzhvDC0h94sisjF5TvY/uOyBlrV491sTs69bFtYRiu/rG+ugw4Owm
G4kbhmfrDuCcUJCseLFp958GVVRqifgM3TaPuqrsILlSRhbKYkPt7xzOW/tZGi9s
34mqPir7CkCi0AqyqfQiChkURkCH2wIITwIrEqac2SArQIt12ddK2scjPOZ4CE0y
pNOnL9rFw9uIIONOJPfCBIgPg/RQk/eG3uaSpUrWQ23ifaVastNTRPGmf98jFvS+
EII8t4lTcMC71FZZDo33FW/FjdrH1UYTYuGBUdaxy6p8iseM5JYaX+qyGbaSjQ0e
2bW7CCXyoQWcSipHa50KWYiEwiFzfoUFq1Fw9XaJIpYA0QPa4YfkeZ5KJ4iYEOIk
ZWBLBalTGXoe+UABiMLTbLce3eGrlYNUD8o+uN6Y9lh4hW17U5KPHA1tQxz//vy1
Vte0r5rEmK0CIARgkzILQIQunoagwIJEXSf4xH2jQ0//MRnet30i0AaFW5yl6A7C
BTt0lUZwkc4ktdY5+pFHaOnRI/fZ2/BOw1HBaJu0c78/lrp2pZB4A1Yts+LA+mNI
yCWWSMZUstxVTJ4bI0JQOeblCE8B91BCbTcp1cBOSRdbjRSWUHmljzJDJMoIVZnw
8VnflEJCuvXQauGrHMXSzofwWignDIMJtdPIQzgrs7r5o8ztb9l2myanW0pSqZ9f
fVms3Y7bPxk8pQz80pA2JvyKo4/1Za290D73611R9ap2KQ0wODtoXvJKZTV8qUxF
jPdga6I8lbnN5GPyQCCBSNMuZJxcV/r+YUcy9XdEeRUjSBsAJGm+VCW/AeIu2Jpc
DPq2VeBliCArT+FUlYiktarWRC2+94Dh29VeNjKxT3H/9gL9GkAeNr1kpA6ZbDw6
BLmviWhCbq6tikz0WpoViXnxjxm0+CaPORzEYaWHjVkUYg15NW9GBZwdeEk+XQ60
4B2Rpcf4K/ak9AMjbByY2vKNmu5+nxpGZW2KGgjTo77fg4gGJgAS8auMCYm8xXho
LYuTljH8b4TYqsOLLuYCsy8GoBe04KeYS0Sdiz0xmc8wCAOdSGScT3jcLEDPd2Ci
Gjbnl30sWmtOqN5AcWuGQ46cVjshJS1J+3FPknJHXYEo+kKKoz2wpaRKu5VlrKYT
qtRUoRIc7HbaeLwXzHRdEHxCZgAn8NGVPUUuzpM4hAvO+ilwM/B7gKb+TmkY7+SC
75+7jF2IBkgxIrDJX79x3V5yPIHxz36hSB1D8Zuu/VyA8lo++PqyswS9fbWmUpwB
6ajuSH+bYQ1lq+LHCPddV6t0pK4gZHoncsAGSOIlBwlbO5Di7oI1ebr+vtikMIkl
AR6SM5zDp9gl3tnt0mXS5nptO7uDvlX5dcC8NFNCYyJfIItEh/5JhzQz7NnsBHUg
4gGdl4/Ksv0EZokXAbptEbk3RFurYTVrmbkGHXf6Q2o+GQAIWCC1C329BuH/Nuvt
Kl5d+wHqXidM7vE7CvQpIN2wrE+FEmbis9qIsE7hxKNGTFmraWlwUXVrRUg3UsSh
8u4Bp05y6bBYcBHCndek6hvLmEGfRG8NXK1M+7H0o4k8baRYH3400sMQY9rvPZTW
Wa9Bhf0kTUQpSJXrXznZqAFsGAcuU7cYK23S4L/I2R4Bk2cJXW+Q+Sf40/EfvpyQ
WZGZDd6rVR5ucL2VtrTBbSijdmYqDiJfa/jBoe1QobVGJlTQME+xrr9mSZuoPW47
eO7auU+i915lvyvw/KKRY0IkNiyVKqx3KY5WTfjaCj+feToxkSMwuCOVVbdLsJiS
/R+BjStAo8mDGI+WVlfXX2fAY58ulwtbmQ52wCL+pmXhFAANqKttBM3oaFr2QFSh
ahiHkja0PKD/e6W5AaC3vwfHUQ0Il1rOX37Gw4JOJVJwtln06g5xK860Jf6naWAh
ZFbNHfOgVubI3Lb/mBNzcNpKIfn/xeTnmxJb2GkpT5xOp65AJG0HDDqpISz5Y6Qn
pMGqr6t/ZMALLR1NV3qEwRFZNLTfkTK5U2GTJSqjvzjoGiYOjuijlAqGw1WLFXgg
SM2kYriMB9XmFY54HakBO5zLPWvVn0F9fytKY5158s4ur3aAXiCxtoQQfPyCZu0k
lRlNbSBhuYYoK+YCSv5yzM4gX8BWyDlpKHfK+ehvlhI9FovvcLgnb4MhDMHi49tM
RiS7bE6dB0nzsx/feMwF0yPbWDrf4uI3UKCntRU9W8omdj44SDqNpCgRMLZCI7jY
g4j7cPO+j5j5i1p6+K4fXhtIkVa/kMRrM5M5mcnaujfpBVk6PB4o8AS2Q6s8pbDY
dOOl/8f2A3uLp3WtJF8YAwCKNwvkgfVPQNzK6pzBNwulJbN8kZhinoHIPwY8S1iK
Q5DAEXAPnRZQNBkmn+GCljV4j0lQb33CvEty66R72UKVS0/VaIcEKiRQXgxGX4Y1
4LHNhBODzX+LQ/7pkBmIytYet2wKEPWd9Spf0LSRILF4X75T0ET6vjV1tIT4zIVn
nDJdSMFQt/0mS8GN95EaRdMC15YL94GKndmPuyfUk85NAuWGt/a4/sCw7IYxWXNf
GW0XSIsQ+TeI8JYxfaVZIlPAFgT3LBP4o996iT0PzfAerpTKotE7wnD0atZ/NpTd
1w1wxUnYFrC6w/Zehvm1c/PrGtu+D5GaSBrtDeebRwkuV0yYw90aKjPMPo86zz+S
K+WqSb7SE3iTAf2TBVZEtz5Ow35ksfMdLAliNudYy/D7PsYB6dNz+I9Q10IW85mN
mkqAOOSf5YOSSHAeuAuiiuHJKCtIa1Oi66H+lNDzdVItPqW5gAilWPmCJj7S3teO
9fQBmTMRttEjy0qx+/xW1s8EA32yrC7wDv+T9TGZeNbd0Djy3T9DTUIc4MIH3AF+
YzfeajtAGaLSWqf0wWJH6OfalIfYfshbgVc+7T9/TvqMfcKCQ7ZBuYrSJot5CHqj
3CkmFp3sTn/lpbmJ1JOkBhe59dM4ruV5j6yBHmQz4jf2bzvxEA3ur9nwRvhDtq6N
IMll3w5N54wXekW41bN9Kwt5LbJmXPMdZ/tz5YOD1WG645JTm2uJf02jPmviObAE
Hig8wPPrDmMRdu1WGy4Pj1FlD5xNP1/2Xf07RbbgMSj86JdL4YzOYaciTvw8EQq0
QIv2fKVN8QOFLycQ9OalMN+41QKX+ucfj1RAg6USSH9/BVO3p5ltYY5x9yCH15Mh
26XXvbdm2Sckya8ZjrNoVKAeJR6ZOrnJAnsMNzQCdDVYMmBSXiDG4WFdr7CG8k1S
ymCOgSo0IMRUwduCBw01+s2SChYnzfpvSTgKPd/2aZDwDZprVUZlHcD2d/Owl7ZO
2mB1o2iqhvteR4am4x6ayBY5dE2q5a7qA6V5TvENjMrvUnbHsAU5YPcLJXnrN4Av
mRNwl6dU9bHhZ58Q6YYSq7BUMX6ZrUxrY4Gpf46khmF5Aa5NP72y4PQc020/70Rx
X9Y1Idc3EojVyBqc7jE66ImzpEXYZmRgTBANQVcRgEsqvF+PwRBgFgf28ND71IHw
o49vG7Dm1IOn6ZfDbnDp9R49pYT4f+L3lOVPGffy8kaQTO874suZqiOoLMDU9ik5
J/jNVwrb79AwWLVLYwSZE1GwDUk45vT43IyYCPJYraYwxCXicNRjr5vAbFQipWnU
jahL2loPat1SdlcJfgGXxRNNiat9aN76rICtcdqCYSIoKOfPLhiJjs+8VVnaPYRf
0XJzRVs1AwwBdnvhzCSVPPBjrXNceoUgmjUxJHSmDirvj/b6E5dh8F8PQnbJW0OW
KP7UG+Ir1P8gNmOrPbNsSkMubI3E8fxMLKcF+THPd9z9q1FIG0PFiomGVZtFhCcs
O8X4IXjlsdI8GrYBDU/dA/FtCF6rx2kbPl2SjJMHUE135wP8uSsxN1LcnE+miE6z
ySz2j2u+4lm/cmKiFHVs45grnlOwCsIfxCfggeJ2UPDjEEHRvgJWVl2EhRPFTIAk
xw981+MNEAwPXHsVmGyU1E26heqsdEESaHyf+InjXn1w6JerNIeMTD+TqPsOqsaF
Jr/p6v61ryaGW4Z8gdxTkdfJ7hqyWcMZl0yy5CLPUkpzVpN/lbbdkDFLnc+xrKlZ
bE1GQPOTv57+sB6dHTHYfh5PfzqmNRl4dmVfhgHeLeOqpwEO30ZuXi5IkUAJr2VC
klnOHg7tzMPAFOuwsE59/YOdOXWKFVt7XyqpZaRP2GP09GjDhEcDo8dcE7KSjjaF
rzIzV1gZ/pPBExoFBOJ/b1EKRqShCVkTF47GEzIT/60mKEHLp+Mi6CNC+c35X2//
G4aFDsc+vorikrsnT6tTXpZoyFid+xJVXbHwwhDpe9cviiJltUaRYA0Icv1VsazI
S696eMltc0JSKMoh4kmhJwBQuZ8d+VvB0avuOYvX7XzI9JEWwL/5r3o/SzWkMMIu
sbCMIoOEUduYjl5Eh/kHLLoJKVkGLb5fRmXXdkvOB93xRF5l0b1WqvIDg3W6kMS0
Md2jwALEUJfy/AdU3wOzqbHqiyVy/b9qlUH1YWdcANaQRPQOQsSiDicC393CidhH
3+UrO8rhfJNdMt9Vbo8PEgzFW/AAB+ZkuK7Ssc+DBH83s+72cK4FW6hgiRFC9hK7
jL5pa35OR21khgjIt/SEqh4HpY2OaX6H0yZAJ6VWQnyG7wny0v9UhjVeijkoLySV
UeHKXlmoFA6bOJKmDERkQSjQGHm4vCmlC4ADGbPqJUZwygsjsPfK1EY9ziRovpQL
EG3DEADysxHCHvH66/rITrcRL9MA74kUJQ9KWpzAmQxAaKvf2O2NGm1iy51YD/Np
8/ZRNzi+oLQ0LEl1ALFTYUe44zayRyb5GNUPWN24IVUPVJuSdoAr/m7p7D5tnvhy
Kp5s7q+FrdguDNz3PvtG/Y9CbXy81OuWqJjXvpjmFdxCAXwhggPYdgJFLMiZxmTZ
2wLXdL+b2DmqBG6KlhjQTxp5vtm4aTwF3DY2vDSqfoTFCoFeLea/Sct6fosMgtqT
O15Bpa0t2HWPaTjeINzj//VGTJJs78HfslQ851oxgPBUeHch0qzX8YYsHc+uIeU1
JWe6OngNSOCyc5F8pHxW16isY2TGc+NtRQOvGo2XJiZceM/76I/bbYxjrGyUElwt
i1uQ40W5TXc2nE0hRogsQuMkpB5pnTxdA5N/D6XZ6xuf2ZpIbzd0YKXfuorGllwz
sqiSTc1TwFpjvY8u82JZU579PryDwwE3wVNDdOC3QE+bKQU0R4W1w6Ktup9KGqT4
fquTPX9p/KNjqMC7K4C1R8tTEMOUsKPCqzcmBz9ujDaCB9Voa1tbtxFU1QAP44Aj
J2O7iWjU4va7MntGcUMY3xU+w9ZIKcUrVL4FH18WjN4+watXGVpMpEjt/k/2VSjx
U2k3PdYucsk9cMlLJEy3H1FasOR8MQmNkoVrLpg7jsSpLMkE/RnoitaCO2kQz+bf
Wt+ZmMEL9gBbVFHU5NYL8Tqo1LxNbJn9Om2AEtvFAqC6pMFUkchmVJGXxRDHOSLG
nlupXt+tLi6aEgr1OdhP1DdcFaWvJcvJgDYIDfyMuJ8TlNUAH5DV1buPneK2PGfV
FE40L3TpuCqdcloBqxjDC3nfvqXL2egQ0gLNlt5qZv4rb51sv2grYCPkgY7KxB89
Gq6el6C8JfaBRzIRXT2vXLknoBNzCxoRAS3LRVtSX7BwG6CtNy5Ln/NJTAGTMg1I
/SiF+gNrlrEAenm6nnBKnEm13BIfa5zPYp/m3GuLZfWmvkIrVRLW+7zW0R1GoOgj
DJ7WJ8OM44WIyymolY4Ai50ot+wtUF+PR9PPKFlqBO1kDf8CVJ0MfK6RdcmjwgjI
81xjUH4sYT8vJmLc9TLCuvQQQEosiMbfEIe+zEhdBfa6R+b5DXtuC3dnJ/uItySG
MJ5D+JDU2pIVRrFgfJnJ5leCTW6Ou1TmOIwNq8vIlbcwVBGx19bYnwGdn0QJpgV4
esJZpguA147THU9Pmgn+XbUv1fuJVhfsqBu5F7Qy01IvTLJWLDFVjpBZqB8e2itq
vT26kFsrWm/VGGxLaqo+jtkXVU2RDZYUWX9R8s7bPIXFXw3X4prII0Bu+o8egmCL
/RXIC4Q4y3vtCkUlLSQ97MPvVIuuzn8OypbTZG3Ud/ZLwBbQlt2mq+FS2KJZmrbe
f6uE+hJnGKK2d0v9eUQeNTKD7/8wfpW81qX7MIvz/56S6NRsQ3q8Ie7Vyzk/KdpQ
0rm4PS8gaoAD1ftTq74sum7LxoOsIWsGblyBcHxdcgzU7KR3xxq/RNARVvBBCQnX
PNJDlwRT0/TgHa5V9dc6j2pqMUzwiWZKc/B4xvJBOEXatla8w35E0gnCoDpNo6Wm
hs14QmZaVE66w3cgdr4Y/exkMk22haLRMiLb+haNzn7V91whaTH6PMLxJV8r0tio
Wne4IrEcgsOhGECrIPOsDfzwKMm1lxw1yCvsiQTu/CGp0Ng4KG2dKYYNa4kCcy5m
tDIFBiHZyAL8QVqB/1Fa6Vdh1sRlTgz+xZE1v/Db3yRaT8Po2WSLtDMOp85uwFJK
AxAQAg4fQgwyOapkygYs5en+jOWRJO3vq82kIIuP3MADWBx4SkETuyv1Fr1htV7N
d+zhWLewSXug+YDuSQoaZLJx1LwiQd8eFcV3Oy5zUQZlzNq3ZSD8A497JoXZWIB7
3tyH+shQO2LvaBPLYD2FPmfBP9lrZicvK/v8iVTNkngFoddnCm+A5bgGxi9ONohR
cO6rGc4BjCyIE95KDVe60bG3LDdaANwHHcEur8hQWwi4T1n6EdGRV7Puptef7H/t
LJkHksfnUzMSwT32LU32WKw3gAH4WOV+EMaofNW1gAnMpQ6QpiFWB28SslSnaB2G
b8l7SgW5hqc/rh4AiV3Ojvo+N+yPKnBc3hDYNPj8JUmOAVOB8/f+r6MyvJBuorI5
69Y5RrBA7kSKLQ4XgrQLnuRLv6KSOYm1rv3APFF7ENb7U5b8qpXB3tbco6qsP4nA
eGVwII4DXdYeemxRtivGxUF99NIMwYUVMrkRqXUl7ntrFwhPzEZvCg1PBk8/MH2J
DdFzKDgjZd6x/vrKoHPqjSF8De1hBI+CEToEW1HhOn7Zt3b98z3hQ+jjT/5R2ARb
H4yxL9SQWB6+4O2YmvQyC1VUwDys105o62+Jet1QzDbPrvTZQjy7R5Jw8m96SoB8
MRZMOWk9t4Qskucmo1oH0r5wJkKCPTbXgbJ/g8ME32xAx6445OSYAwYBR3rZHkKj
ol7s0kW8SU6Ak13R8bfBxNMkv0Zi6EI4+BZPWtQGduZLoMy2LgRZ6JbAtulnlK5P
Upk5P48r0YQfikfVMdiS/teAnBxtdBI1jlm2hmOfMvUNnM6IH5RE3XrsH8tNugsb
RjTLOV04P+DFla1FaoLI3p5H3om1HyNVeLnAWS8kp/GHLWQWRbt4WqSCQeHyzxS4
CP4ilJFczmThiH8TrjYbXgiOYbVspgw6unqbxbgQmUy40zjwdBgv2yusRD63JTRm
A6cEX/jIxITxTx0Ooz7H3hM6s0hDQrV68yPvROUPzduULjUaDiW/ZJdjRbVWYQ+Z
4NbBGiwJaQtAgp8LMa1PHB5X+X5k9/nW0wYXlpdc8eHxjoJvLefZUCG5DUahIS9M
81R42dgVjfu0Oy07KqZ4i62PzlMs79AmgT/8x9q9a+/PotApEUW1ntZLdOVHJbHJ
bpjQLWmjkkl/Vslm4/A192nDhMqqB+yW8jalEUYARLaGLym6pDDSz8R7FYzB7BYG
UrrKhIenQkbmxn1CSAwcbRpWI/OatK3CBoVYPUntrbY63IfS5kVzyK6O0YlwlMnd
0dDqtqYmhiHspjANPcIcuH+x1Z80fExX2x4SetOA9h1trlvMsZdg1ckW9wRgmBwB
TuYOQkG4JUg6USUbNE9nFR1lhH8bqy2zfwtxPomuJCftRyQnKi5A0eBcwSZfPq6M
9kznnrh9vdF9nwi0qdwVgROiGypMq8hDvN5+keZhLziwLLAfM6CNs52GlpJ97gG1
GhptJ9d+wgyHVvqj9ecHJlPeOu4dBfrRi3tgZqosM9Y/SatMIZR/NT+MHcoLlFDs
qSdEbgD99Yu6cHf10780hAmesb9vknrsxj1IyW2akllrqqDiYIMXfkpMzSVnKNW0
h5PIIeESLqft0RYmw0WOLBJvuwRtQpWdLrG+6LQ/4N+ggfHvGK8e6FoWUFessMK7
hsP/4LE0eqnl85gpN+2uXsDJjhyTSCdY8ncTCCRtGEbQ3ffKxHyMVqrPRGt4YFMi
n+UV4CBVvSAaXoz7KXmeE9xxRr9cNrz4rzZNTa6K45dr7nKEkTpO3yqABkj0l5yr
IJasY23X+82MWTMh89gPmrmnlcrSHl4wvpmjORzr3HZeUkUS42WlJEPSqCaBWOiz
MSJbJkjfa2NTVEvsELa116VURvW9lKr8l5Vux434jcMW8s5IOaEVqCujhTw3c707
OWewwbK9sjNOYejYiJ5w5L4MD6bROtjxA7j2f9niQvQiWcdV+0L8+Fq5EbWhL8v3
++NfNFHe9lHvnvyrH2R+gtOwEXZ/qGiWptllTHndFy64qePWYJMoek/Ek9vs0pAy
NoAO+n9pXsruPLKa/+tgorH9eHTuIOvT5ZeMjpsA+lzXWM3ifQwlpH+dgFKCZmvW
hw8HxmqLFntuWeq39tZIvHsRlbn76bH+VqioWfLYAeTEXh5HaHWcSw66MTV8zw9u
+6nxftmxPqHJlnqF15hneMmkYJK/2k/DRm9fOIEsccXqEnVSH18aQJUuDBlLNw/1
H3XAz5KZutHVqullGj0/7BtMdmLIKjupriRwdVGluuvhe4yK/amvlo8vPcilwzWS
pfCMhoIX1T3yMWtpwyvCAsSMGtNArSpicpzGBmBac+QwZgM/C4fwFQeHdEGmIEDL
Tjggz4purQ9FJw18EGi13LCridNfkBDjzQSqvxkBV2xEJxZs1VlVdrEMXu+clCAT
f/SCFgd/rgNjIi7YIq0/wEXNNLeTOmchiueYQWey4jpjPdYjc5T/Q2bm4/I5/V28
4tHX/+dnzjMa/WRv+bftJlbm7YPmWEju9gSJnOMfb8SZ+Sa9zBEIVJgXkUcrg2KC
Gh2OqkCkPqMcFyoUHEUNsX+ETim7CP+2pUWOyA7rFYt1wr/3p6Cxu7vsDUWrUGWs
RhdgwNKT7CiMOjCMPFpvYRtBktTV7o7f1RkC1z/CE8T77vV48AyeVviDY/PapuG5
tW4S2Z0/71Z9U7DKeYV0c3AsemVuXcO4UB0YpEB31D79wvveQ8++IjzCOQ+78Y59
9G4T/EJnzw9rN8znauocq26/C45grKD7jTco72dxIMUoHi0CaH3tWG5jB0IR0N3E
STKNUmdiDbOmSnpX3qY/bNzwa71ncaORSrEkHAmIV0xQILfRCvwoWGXzr3rYScNK
NDgc+1871l9eEjNRwfBFSdBe0Q8JnKIS92k2YdtCz3m4E+27b6diEQgXwBK0qRcM
IJfNmjuzOn7IMQlkZkvTfxYawuZTfjzxWuQZPJU3CnPFPh2nESVqfGyO/ZCpOuqH
cwvgcQ3eAp6qupfHDpB9uLeiJhfd+JXZmYV01ixEMjCI7dGw0SQcWMGnOu+mtb96
esZiSgLjv1dxLaYtRrx1DIQ3B8Ln/B7W42Z3JhfSX+0FX4kd9FphWulZCOCWjSbE
Po1fYWOdUwhK9Jz4XUfJiXjGwuSKG9mj5JFVRyCsw6yN+tvryiJUJnaRaeVZVxV8
h92ftf7/ZYtlpl20yV6jNIoawBQtn9XOC2unpfuiwIub1LysYDplFUuUnxOuTwty
pedbXXL+DpSLXnkpaNaYFz/kBuLSOyEvsf+8Bo/sXVYk8ABKPAMhs3WqNNFzbmkA
sqZ83cANmc+OWwFBcmudlsosi668smDJTqzxycqoqO0X+d1rfWZpsak2hHJvwx2/
vY5napm+rhRNAOBOA9zf2ZuEkjN38fGjBMEg58+BWr+EuqvI4hC+0S/kGxmMRMZm
X4iWiRkIqRq7Pye5IPQKOPVnFdJIl5auZTJklvwGScF16ljSGQvHgg+bz5SKuvss
aMaKVYkmXYrtsSGRtwe/vTlmkE7AocscMsro0+0EQrDbPOnG0Gg7jVFT8GM2FdMx
K6ZgrlCWXiKUkdxrxCXM+Nl/AMhI6MvZfbY7e87pMzM6YSYWFYfdSAjJrq5u9pnJ
5CiUKG0cIhPsIMr8wH97rsIlRvOibCFSJwC9APbnvSrnGdj0PqmWfwuENrtizGqF
9YByuTZCQ/GBWJTWg5aeGcPRSKtNR0yfPZWIsh5PYkHD+pZHs9tdGp1WAhhCUwDl
zzouPPmki8bEmxomyGZMppAdjL4sxrj4YIH66B94g5+4pPoEmc8B30ZSn07sXTuH
SFkAopzzZ3nBMCMgYxqGlHuRNcI9aUQxXWHdcBSOgWzQssR7i1bYVKFQHSMPUpW0
eoA9P52iw+iIKBp/zOeW2wZUSjaYhtYHSJQk5QXtfj8z9lxkHqrO8t8mWLy0M2q/
lwe/3cDO8FnYb3srMlkDI79htl4m4vDGKLqGBk21DO+NRPdEZ85hsnQshAfp7S1O
G1MBrFSdk3Slohg9C99MOvC/9aqpMY2ahX+UNxCjeF9luNDiyHI1rdFS93FYU2rq
rE+YnNdNtvjbW4YnYBP022RMnKHzddIga7gvGMoK7F0XE9sVrvXqcRA2uMHnUXNw
9MOuCiNZBXAiI72NOHGoKBgFYj5ChPSl1QnVENOFnursh7E/1CBJKO3x4guQzvyJ
lCU0gR+5haREh2pzO56Kf9ZsZv1empYDpMJSfHuIxepPYASCoeuZ5Gu2wEpI6MT5
nfYqJSYNH6VyAWq1kKxGoZ6A1L4BmluGrKYMWQ6M6I8r9iQoLuuAak95LZMjPX6h
3Qg+C/NIhhT8ABeRMo6XcCBZpGZBmIfbmw/1c+HRbsJWwu4vh3z1NMK7P/M5X0LA
4o3VKX7zJ6oW4ErzM0FbO83VB76KLN8qxLnCmb3hK+rlqByNvAqgdcvH4HncAK28
KYK5GQy/BGvaYbJMckjfT4bafPSQxVrHoOIQUH2yjAXdTCk9rHG11TQg1NFWyUI8
iSWlCNVoVwXSp4SAA1F+Iqw1io0vb/T2lNvvwYGc0VkhGuiRy3DXVNZ0IgOIvEAH
vj935uRut2KkYHlUhjqPZ0o70UkmGjGy8I58OJYBudeNLYJ8UxES68ns41y9gi9t
Rp6Z0y23nQBOeoVOHhFlQRRuoYmlSqXeyGG5T4iV9lJHFxcmf2vjc/Kn8wmZld0d
7sE+Z1vkvO1q+lJaWKUJB31qnroGYkrsefCogWvL3LZh56IVwKg7T+Xmu1rfV/Wh
ph3++RQIFK8LvREosP9z3WLG0JMk93WeqJYupQEKl15gbdmI2XmwMcBElsS5kwA3
LT3EHcefc/KbfK6RufIXdiadZTYEMiDWj0rerI3OO/ZHZp4VovEkv4rr8Sdx4jPr
U8x/I3PVVO5UTz05KbsFrcn8iPcfLtfqi47LTg2BSZlpoHyIJOPe+KW5tmFktbzQ
+hpSx+jme+IbRpn9kjGOD4PcjMa/7NE2a5xGAQLvOzLGw0FNm615Hc3xF9HiuM12
404QvPozbd4oJ6InqYD7SIQnMTiwrKFxV0w/Oescy/8HJFuJbylsWZ4+pNpuB8+6
XaLkPDSFYUSEgDuBL2w9mTYdbJUGT0wgFstPY1vcNZNJO+IXHAhLovdbKFfpIJPA
fbTKj20Abs6MXJnyIfemCrjHwJi0Af5LKhYm1f/hTR8L2NfkM7VemtZHzFJ4MW74
x3HJGz2ykt6C3T5XKSDNxYoVGN1INvEVks9+LdBxNYLmItNbFXRuBauVX9VrO5RR
pOocVSv6v7+0+g1wPH823E1DcBG1eNxZgWxu6Ch6WsErI0p0K1xWxmapbvudAcj+
DOe40iMdim2Bvyz1DH1fJVyzLc7f4SA6byjrdZECIxgMXWYWBelhEOw04/FmBxyw
ttsbONN51n/YoZLIPzz7SoF3J4pACHE7mmkIuaaf23nr7jjq42SiGUJoRl1+qUY1
dQ0ivIofzbT4Gfu1cPJ2ybYPutmdFSO7G7KrZLfo6C2uozAX+hgxkTalPANEDAxT
UuE2PCupvikG6QGe9Wi4uHQdpN8R2oX8Ux8XGF3w+kub1+Pwz90GWmOE+XWw6BTS
YXFVF1rPSSBlAYm+a3NN3Ohn9NQoyk+7Y9IhnqB6bfRUryiJzaVqBsj442Kf/1YR
xDDafLfj7kILaa7a86kGiEBKP6iWv2XYCBRm/yZ5gePQaS+XUp7GZda6K4Phyr8M
46fe+Mp1APtXF5UyMg9vXEODtmQOwp5tQUaonpns0SkD8QogRIzz1w0IiU2AIieJ
cFOevivm8qpSw4EW9B30AAJMl6P3MAu8Ezl+6IfVmG5LkKV7d85ZgY8JA17OV7s6
T3C4yq8GZsd67mXSyiSQEQkieCMPL+bSsC+oipL6Ae33Cd/o+gnFhejh8apwgftM
vIHQnP3R6AseM2OMGD6o8n8iW9iB4hndGe51loyRWfAe7yEpns2vR/2MaztctW6C
NZAVPiaQaO/BMM1X8sNg+KixZQU+nL7LRQnrq3w7h8lN0Dt0TDXUYIuYDGR6xiOF
gre/r4CJUBF8rgHWo3IvH/LhbqW6cpv+IJrr/Y8DVZsL2XH6ApOxvw3Y4/PwW80W
JA2FZBYSGX6REqOL5bbHJjKhp7zF6mlkPNv1rYgyZbkf4IYc8Hnbh0RCFIMXlmpp
SWHTo7z5JWvnSxqov5u46zeH+2S/Li4OG/7hEXpDRbg0yg6gXMbPMKfSO/BwVzxA
jKyW5bwpQ1YM3VV/BBUTI6iJfZ/umXKJqD6Nab1g01YuSbKBytRZzJ0Ic7WbFHu9
l0UmY5ixkvH5rScAswYFgHWFl4ya6aoj9EZXSqrXFtZuV/XnHrq5lP7exBCf7Xnm
3NJwqdxrmta0Z04BVnXDAkDvKWVSlfLOZyhKfXyCE59MAR5T5UrbRR5+cXW0Zal0
i6qke+dGFv6bNSU4mDoy/A/DRJat6gqaQ6K1I54v7xotACIxkkoNpCCNJ12ZqVkn
s1xKG2hx6Bp2IrWhVopOM2PLIaXktKwV6Vev7tSwonyVDMim2NoShUjJQtzdW+vz
0Eu/GYlVyeF0Vq0rJ3JapOjNncv7jYSut5ZymZ61i0eE+2gIX58OkRoE+3XMztJo
QAzeGmoL9xzzKt3piJ9iuMzYLDasqludMK47b9JRR6mVjysLObkgMqDxqNDyFvkf
ehoZqUuUXumPRkDHNjY3fISoeTizSO6Asd9H9mwfBLPWFY4Z5K8H+4MdsZeBdkYB
oMWfDsIS/2Vk2E5CD7GQBSWtgg6O9EjAaAmsts5dodwUe9bjNXDy0IjZnqW0go1v
BamclEYkVxmCkaEzxPhO0Ogl+TluLEXcqBMYIC2pOxozR1GUj/IZ9vvtZRjbym0v
eaHm4eQ708q8ow7vcVb9SU7Rvg8WpvdhLPlNSR3q3lIy2dtdAT+89gVQjLAL81B+
wuXUFv7BA9Hd3pBvDqE46/BcRkSJzM8+F4CvgLF6S8ySlLDtYPUG2wNN8wMPwgyO
zeBvX4T+P1vm5X949+R2iymdAaFYlAxzz4Te4OS7Rop9J8NLQfyHwe3wZDKKvUEe
MBmqFC+x6Xh2JJ8YvyBYNz0Rmtn6C7nu8P6jwENTBcqJMcZ51SH7glKrfVz0tA78
+KxefMQ0lUy5K2brPqx221QFsbU5Km3CZY2TGcsiNH7VQ1guEMpMCi0Cc/Uhs5Sr
GG4oqTJbaPVNj9YiBec4H07vkqRyK188vchc4Y7bU1HXvTdVt6fRSE7BsyRHs84O
Zuq38ClffsrkVYxrj3kMH9/IBIF/qryeNuX9Add44fAQ0KuZwvxb/85u2lx9YNoY
NahJz6qRSHOLxcVO1l2RKuIv+R3bGwfAZkIVo3KZicAhaHUQYsLS589Z7bOdsOWr
6T7bIbCOWu4zulZ8bAWNz6QjcMVxCL4ZqoygPvYOHV08NZEYT4N7Z36U+zt4o4W8
tB6olFnQAO5xj1fUeBYboVjX+a7Kuc5tIsvnU1pQZ5yLG7DyqXzZy59lW5BmVflc
JlgbiMz0yQWXJc6WKhweayTd6VWWe+j6fW+piEHRtyv7x/WSRuPXbIsGVJwmePud
sm1XZpFQ1RBpqeeJQ7tOQ03SQjp4ORvLl/b0d8f961vM2kZF5yjMvRBSbowN79bT
nL2ApyZlZjjTVTU3h7sd5ab/sLiBqrwrNvmuCisf68FUN6ApKGUoLYyESrG8kbw8
McripZ2G06xNsluw5LZIpzXYZBX9z21T3bHOPw0Q8TZQsx++w2L7liuBYOFFkrF0
WWFNR9TZWMTqNnrmO24mpy1USDVIoVAxZaVtUaohvvYWCIyWta7c48i5uMI5xiMj
jNCXye82BhiFZzCmyjbswKaMXAQCOKQVXjpKZiBaga+hEdOcYUHWWbN+GImQ3Uhn
DI3lo8jsP171mstSVI1bNv+I7JNF6At5WFCSPWVWsWz50Y389GH1prXN7ZInNC2P
Vim9bLoVM+Y9Vj7b2LcpHysktM38OwqxrinNorhQ9dnTPMOFSQA11Vxhp+CnqjG8
FbuKoJGlK1Fbk9qqmtyd5/TL4jB5yWS7Zir2eme5PfTd6lmWT/EFsOZacAYjofL0
QEy+B+oxUhpPZwFdEOFMBqY4J0rNmykTolrWBv1q4k282Bq7MZvEr3UeTQd0qPZs
7mI4jlkiANxSADr9yxkzeBmXuO0AtabcuqJW8mTP2x6vPJaDxRSpfnjKMzyTilJp
vyIaw0UY04AtKKW/djv/5QkzKlXk0fVS3nnJYDy+SALIaxWpqsSnmImxCCLALmqf
+SDg8OWxxGCLTYXy4B9sx+GRTgBn6b9qFYB9hqHWNITsyCA/Ovy7SJcQSt9bjBjc
/6AK8Y+L+R24q8uytI9CuDU5yBSa4O0nvkRI465c/pV3lrdHjIIp6GotzHECXuRk
AG35BifiP06EzjBAFnJOgVrQIimnRANoxR2DFEg1DDU+NGNioctFfdCBotHpfNsc
AMpEBOCKuAFBnkCL9wGwaTm8k/a7rTcB5vUVbPJz76d7y+ytQr2rCSQJqbVD3Qjj
h4TlnY4p/aN3RNhT5mFsw0AqZROVCDf9ZaxFfMBCQL0aPdKz1uc0yKMJgrUsEcZY
1RVycoIexBHHdb2cwQFMCZs/oK8OWGOma7kwDIsydzcDqk1oguC+8nVyIaOvVd7a
amHzDNYlWxLe+0lKUIWt8UbDyUV/osB9VHyytdMhORDsffDJnCgbEmS0RdwryIGL
TX/O+lMJRecj2xb+IGthAMdZSuq30AZVgKAQtL7CtLqkZbdVcwH4T7+undK9ZATS
/yfZol5gm7SIpaUvLqhbSLwlqmiq9CelNDCz5yeb534Pa2pTlHPDcrZonhmcpQM0
PKvKDjyoUXdd2wsv1KN9+WUUUBe33pnpkS3JIH9/0zQJK6vOANobVdD5fSDKau50
nmOIVbuyzMY5DILAUneNkSpecszY2RoamJY6fUOF2hRbOwlQkWDjhsL/THWklK4p
e3LX5KSgd6JeVjahq4XW5Qqjt+muC+dcVQAAe6SiYTEHF/nLgYXLYFq5zGO7R5oA
THADk/ZTIy+8q/nVoc3IWxk0H/Q89Dv9INr79HRvDqhPr5zhZNxWD/sCBB7zXXUr
WW4j6DIhXNvRlz9dZQCKC11TmjnHcW+tfOhaYXyUt4axUi1NxgsN4+beTyBnP5zx
gioV6GnDwPWNoF/U4TMm30w0mOam456IRaaB2ICWN4QJgBeuwasQO0hgbwk2d8Ut
jO8exLPVTADkQr9koE/GnUW91UX2m67b41MQjqaaXU8dJr1ByqlFAAbPP64HykFA
CNNlgADOa2GC2E+wCfvyrz4PCCkJjBMgvXRJQaP4G44hY/GvGnWnQ0/2zCFCVbg/
9qly6+1wnq/mkdMIdFTUrMxP537ke9QzEet+xERwnaAG/B9b9ETSHAqUkIwZKS4v
4ff7ayBAHFI3PVjI0kZzvoJYBJECvLGjYRk7JHiHHDMKA0poE382mrW9vo485pUG
u1IsSJAGO09Ym9RixYh+qUh9tmYrlA3+JHD4iaHxNkfXdnNKGabEMGNgFXvwLMWP
hWcgxFZ58Qxk5gfdSFwimAeNHN3g0Ohm/t4qjHcfEDnsy9jLM323Vb9b4LGlgMg6
qlUwTIHUfUeLuvWRROi7fYGufJb30d5Io7xhNhUlIR0ZapJqkFlZEeNuu+prbpAI
RhAVtsqv977RNVWrYHNNiA9eVUY8JpNeHBFPNHQJJykX5i6CFQpNbjdqrUwYRZul
LwYurCZuOFG6uMwkVwXyBHizOLfRPMdh9vG1fucLidDtPed9cj1BOGZJs07i5vD5
ZgXfAm3U/EGqUG0jdzjFOJ9lqAEAUb1W1IZQfq+rx6PoBfhswAmH8ojld6bkkt8e
vl476L0r2G9EE7P+Bvns+u+UauOSRyuse1kamAp5n9KBcElB0AtKAllGBPOChNyy
lbajGxVcshtXY40JuUETRM9TT+dL7/O8xuNViRh9KhhF38R8mb1aI7qVxUaDSGPz
uk3b+OYVY6NmYkofZjWwmYrBh8SHlevFjmw5oTDkd9C6Kepjey0HPbO6BkJlzxdP
9iCDNPKFrlTy9YdneV61oSMNblKdyM3Mbj3PS4+KOhXKNpO6bk1+VW1P4zVpZKvM
He8c6A+3CrXrbGZYjmCXA+AO4t01911Z+UUWjkHQZvHaMpWddWYzKugrqsfOTrgI
cvGffDX79u0HuS357L0qff62va1BOxWI+edx2ieVgK3eDSdN5ArARRCT/kmSNasA
eVac3X8zQY6EPiW7ToHOUs+i6F5cZ5koBfQ3SdEOguXDDbaVOInXCP8MhTo+7ywX
7Rg7dYfNNvidNbdBTgmGv/fF3Oz5+Nnpg2SPWb6/ub/Rlwq5Fs0sE589k9gpvvpW
QrlKFJ3xx6MlehOqiTr4aeEhW5MMa3VvKBnITSawiX3P0QlgWjgeR1dZ7SBEE4Hn
lBWLKJVegqf+KQfsEIvsmLnnWbMv59rm+qxFi46Gz+zIk6OFkj1RRMEQfOEAMxUD
zossjOCmyY1RNXouw0+56qtO2q6CeZq/thOYfySEosI=
`pragma protect end_protected
