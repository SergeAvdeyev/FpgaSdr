-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
b9UCNOwzWB/Utg8EPflypX5TR2HlDCVVybdRG3nmqaL7VGj44znL/SI8cfckVczDvYRj1r/e1j1j
fYsG4kfZQR2YEzoMjbym1ATdNGvbGWGkwqwR5mPSfgAMnjboBnR4fgX7BGLvAxSJIoR02a2f6EsV
jcw7EGd0cRNIQPpQc5Jf4AI528KmjkPAPKN3Skt3CTfdsrMZLtFSmiJCF/nZ9y2U49bNgpsccD8A
X/WlOTY5jIhVkuVxSntS5DiXaSzqhp3tPRpX1b1c/h4mn92mt+0cebXZoxbROoHHK0DR6yCijon6
h6SWWd6zBDBQruvgc57m20KPUtSEZrWyZguA/w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
T9d79fQuvKors5b9Or72e4M8CQMIrO5Z8JpXRY0qrHgrrYE7THAg2oFc3UJTBYEjVpLwgF+CtS4+
Gmn3oadd1Er5bWelN9bGQ4XMwbUNWezOpnqiCnXjh5uKvTV8o7NgIPcxvgg52daHJK9XCMJwn1Qv
qCXeXfJaUGGNMlAp6R+jlz4ckVoiHgB449OmZMHnvxCQZfiIM81LNBDsWjCNh8Di32HRuozJEcAe
svFvoqaeukrv+gff+OekaX/qO0HC+yuxxL0a0nXcdC/1N3h03Tj4qlZRHEyHhMymvS8RMKXThz2u
E8ip7Picw7BOQzu50nXQku4llMSquMFWgYgF77koUR81k6UiG6xnHRNZqLkRFgTgPGWyOLhgW4iZ
eyFahb4ZA+pL87nqdhivZpRb6ngRgUC6dhya9ZWMYsHVYtukTm3qOgtclyMuT6A0MafhDggudKMU
SxSTbjrymeq/1pBVDr4pJkXw1DRfz1zOxAyMX+9RPXD9VyINVX9AS4T8jyfMhIbVjxHZErfbu/Px
hXDk4RobKpQSyPCa8/WZzmtjammwkuWyxHSQfDg0mLGEaJLJdCuHCdf6sFR5scRXWllTMB1F0Fmu
kKkxmUO6YHRLdEo8aDeKOyzOWOLQWDCqj6qEn0LUBSqIapiV8XoUzZj5Qj+T+WMP9AFmJ91LMA8b
rWG3FqBwMPUWr6NO6dcvRpQHq4CBLf5YAF+s2j6s/5CfPISEYvBlKwPh27+5DDg1Hpu1pJR7Tf/6
tZD6reaJCKIpQJZw1x7n5rXGEhHnKS15+6KM4k5t7eUk6nSXR/lqay6atJfL2F7k0kCgWZ59CU+k
9fBpye+gr0iPqG1T+6JueCIwAxGxyMowqg7I8Hau+wUZStaUsE+IgNTt5UBab8EpBu/uAaKymNMd
vKivr6lrgU4UCtZIriftFWJyxigNOJ79vBqT05H+htjLCt1sXS75XS5SWDk2ivhfOkm5rwRPMrhc
ln9or1M4EDSvAN5XXrDDUizwm2AKyNOoaxlAWKdcc5FXa/YvhqQQSZIWK03WaPo5iIOd7zR6e1TD
aEwQ0Bn/cP7t/oVDxjUJGhjCeXT0kf75ah64Bnha4DdaYcKa32tRWbOqRGG2459vZYlfTClg7WuW
TDxE6x9elKwrptMA2zDe+pS/pT3R7iQfigSqw3SElq+GXH4Oh8DjMIjqZNapQAOtqeIioZpNOUwz
fM+aI6nipcWBpPb6mpMw/LyphaGSzvbDK4D4Vrj9o3o8fEEBCcYL0sjGHmP+R1kPXIsMmWztH3uG
QnWTSfzSo28OEoucC4SIFU2hbiGFZPKCKf30w14yVdHrNL3LtAN5RLzAfCA1CkCGqVXsvT40eSLb
96mZxvfWrCKYhHAeSWlUoKzpY22hKsJEpSRSqRzwTKk5N3X77XhmzVs5Tc2g1VBlh52keNdL8EYI
fyuggi4MLC39GmYKUHjzvZpGGvXPe1B8sU3JqEk23SJUNABzWYBbfxsHOP6G5DJE65bi5Uzcwu6z
nLYbsQk4hCszEfHrPRE3iWQWMUQ3JyF7s4URV+gxKYB1HyGiwASzpIpBbSeSOjt4wei3+fEh6wY0
CPNrgar49wd4BJmjfTVfzCPMS69TZenUhAO5r5Ltf/+QjLBjMZUnQ95S2wSJA3CcSO3Mv6GdvgcZ
tMwZG4SiF+ZU31kZWvNhOvCLWpMptfLPeModwf4cO6TrAm+kG1A6EK75Pa3mR6CH34rtX5FTRtP4
uUBEP4k0B/uRRfohnk1MWPEySeCGo50AfFznPjeQh3dLoKDtF1U7jNRmb1THYVLSA7SkZP09Xgf9
r8VEBrt16JzLztmb7qDRVPidRueyAx4c3LLsaUq7g/2j3uQU5k9riPzIb9H3LuQOXVaYRNYkduga
YMeMyzK0yoGrfa9ac5aFTRuwS/O2g2iZq4adUHfkEaR6F6G3myCBH5gXv9FyhxQcc5kccyNxUj5l
uk3DFEOUIO7jXl4/S73mYLNzpIqHbD42N5PKEt9DEAiF+WLdqMQv/J5aNaGN1xnOElXb+0Bx5Qw7
bQc+ekEoJpJayyK4VWcIAD7BzKKsasS9GNjO9nB42R8e+atb1QmIWFS0kq9d9XVyU+/CrkDFHJCx
139GZ9MWCvUp0C1UwXCUYK8BDerbZZNTE0hCDoeF5j5KG5XUZDNCeWlzFXUfOHScF0EEXSAEigO5
k7mdQFzVN+9RR0zJNxBtNHMCEz4/51hDjO6VIRBM8OJ/r2g3bDP5IN0YhNEXrFT1gS5BDZejC17L
AMtzi6NMp+99uc29uHFhOmst3DjfngOrGUJ1Umnquz0Oze4YS5h4z7OhrDsxLnh+gKPbYnzFZmrB
7LxT/Tcbl53DxpDH87H5FxChc/PmIT0JZjKQu0EvJ1EsILQblBx+qGJFUsIOc6QdSnmLrpiU2ojp
8r8vCoISOsRcZstprtwAnjWlseSS+L3Y7jAw7qGNWNCztmcl1T2yWmUbsP2lIOjf/jal90fvR3ZG
uosIaBIPvHMKam5DQztNepsesCjkCSUCFpwGwjFUekSDsNugqLX+jgslRNby7UUnvpm4Et28+q4N
IXHb0eK2oCcxxjkAha5615ENw636e6wvpyVpMhWLSILvey0NQ9ONBbutpmHpcFdRPTMKIMrY6tch
9Ly178ivkHCVCuwIFDSejsvR8LO7fLPf10QYPPKSCatB6ExwVxhTETAemY6i+GmsJ5PAo67FV6/K
gQxKODnjMyUZBAaSyz58Gwf0o+W5HTin/3g2+5k/F5KmB9GUORMwactX6IxZEp2qTm0y3WrRBMnS
2pKWGlleymaiQyX45Jv51qQ7V7fNL9yk64x42XBBXQq2TTF+757PCXx9zph02zu/gN/JM7WF7ZRe
arMoxkU/llcS7BECCidGTO6yAwN1Zkuzkq7KRbGVZRIrgUgMsZFgZeFQvE8jm0AN7ZaVBN9eLwXy
RJIX+5QfqcRBfB0f7jAQEMXOGUaDjTewjOHQ9Y9x9fMRb4eklDc3PrEtF2vzRpR2NNuk8VQRt1an
LRiLDRfQ6+wOaEbkYIVJN+hvISslldxi+aOOS7f9KYYVhgu6BC2CLP+cm3Z9U19iR8RvDNSTek17
1qw3Q7fweSsnXbD/rva1sfC16lf+T4YWsSrTDhh06G3AxedSPCeLyHpRzSomZpamuCmpN+Ck4y6J
KyLPlv+KDcHigZJZKgugtZqLn6Qb/QwSLh6cZjnWWZ+/4G605JDZrDnXHy4rxdGT0EclYwSElwED
y9j0PE7x2tatN/1KoZCle+kWWPXPLrEHLpeptSAUPbxArravhE+NnoZq9xHZnnjKliKcW8GRcIDS
s9r458UEXMNOIyoZNrLoNkTSF4Km5LQ3tVEr3fxBEupJNnEW5NevZknVCJYT4hQANPkx58mOfR1v
cHVVR0rLcCRffb7R881ILHtI/hQjWpAtB9PI/zuweByPBo3DulsefTqVzVtWNcK5VRPwD56pnl/S
p2LPc2zdsMvBrSrRdRrDCIZ4fmgg7vywUZDd7oxrHyhrVtHNGiz8DDg1RTQ69B1h292NSduYS0U3
AbHeT2xuqw42l5YHy4pXxt9cDR7oNj+S1vdsW39Rk+CRb3ndvz08Pm9ybDESqRS4F9y5gnwz4ZMi
5iTKXIaj4a5Xs0ZLzVn8l6PcjPEkCMLYH65vVYknwVKW5mL70NiXJVdkBDrzsRo/2r+ARAsIaMFP
FPk4imRzLwXeW33Lg621fNczAzzgC73pEACxzLIvqNM5W1LWZ90/riW1AYwuW5M8PfT0vWpNYrZZ
IG+EED0W9RMEE/bDNxwr+5AZuGb6meouKQvYcNVP1XR3I3ZUIqJz4B6ezMuXUJfHh6ONrwJ96gMT
T2JdUHnEkiIaakoTZwLQHR+Lwoqfd8yJTjxJypGRkTcBBZWKgnn/juSiJJV9BdMeDAm26S1/wQWG
rY1VtZKhoULLdu3GSHPhgk1Hu3Wtux7lhvUxy/OKC7HRU7dl6nT4dPTiY+L8qMOSp/FSqzs/r+ZB
HAp+q9kbdXB46384rsXUtBfqzf76bPrJDAe1zkuv0xgXJhNbyYOHakTbLBwQve5L79cJz8bC3ZRQ
auL+n8XKtiOcuglEYQOSnnGUUvDUuBRUXpniNXwLSvXVRlr1P/xXj0Vm+8nJvI8zJTRoS+KSec9n
UHX4T/dwpTx9M3aI5LQ8PqvoxGfHh4sPacGDMGYqMIxp+lm5xRPbvfbwCy51kJBMSi5q1rQZNHFZ
wOKNvl3OLxmi7c54AoNjUi2nuPQmgN1BHCsiE+RkwmYz79Kmy+rcVsFoGlj8nZQTaZT0ejwYAjIF
cdxGaJkCPAye/uSG1nWHr1IlYmHDI/qB2RdpvmdprsFG8hA8HsdVDbSdFPXN5imK9D7Wklnl13ES
RlXCJ+N7wD2kXVPKtvLv1O59rg+jOOGATRUinvzOn0drBmJGaOhM3mAuAowL4e9I9jU4IqLZgs0H
MyGDacYPYslFz/WCNxsWA5clGWjMPi+MgJcI/3Pc/nfQJumMupPjibaJpCkthCbkVxKKuBh3UMCg
jWQBhVzJo/md03gvgwfOnxKk1CvocG3+6XcJdKw4j/m+QFad90rkkjNinS0idFB7RJ8CvD7/hF6n
JEtGx2MUmBz6CzT3yBwfcYTvunHhRwFp31u2qQdp5hOFICNGbacRI0omNXR8CX3nyjSl5pAvtrjO
+3sNVeSqyswXLDTg5EVFNh57uvZJ30OqErS0LLWqjtBu0s/QLBa9KMsvj+DtYgvz7HNRyKn5Cm49
iCFI9xVRS3UNd3Dd9AvP2o2ta0VmhxI/Ws+ztlmVrABStJa0tUIDXqmjjZwJViDhygMWAJTF1+S6
qoBO+8lrxbhdh/iQ4NKqJOsftImctiN1k+0zzO6+bSHtwu4+eNPGsFBmlG+k7VOQo0TZx2gTHAG4
uOMcULDIvHmiBIv669R6Nmg58Yp38DcGGEwhnZhsXxBgZDCEWKlP23awvsLtICLZIdLoFhPJpS1O
ejzynhEKYlumgyw5I5pLb1DKKqluxkP3ZrRECZWZ5Db7wlvSstAwH1nVpcUw19kWxZ/K3I2KBN+R
4VhybA/b0k2M75BHXyS21/SthA7p2Z9QAXcZRs6AC6kUJpBuGFKp1sxudRJrRz+CB9uEchPBuhXl
6j7Jq7iY477X+yuOg7kkyMRy3VTclxzbsS17gSZVc3quLBdWj7hS0I9Mkc/IAWLMY/vyQC5gA9sp
uzc7XUk5j+qmartYO3Crx8XGfYZ8o2siH5dcmzX2G1zf3A0nHsTs1wcffSidj5gouSIX+hmuGbvC
ITWfWm4hVo+FYSslaF9toYD31/08sYU4e8D5ICknENTzuTBA/NqB1+TS/O67rtK4SAMjNA4q6TA7
4w++8RdA09X8oOQjT+bNoYNHnR2vUAn/Zqp21RgZfVvWZb2bHvaF9fXXfz/N2wyzsXlIheUGDMfl
ClguIS/qmAASU+I57cyhXuhLylgXdit7ewghfGCnoB0fku5AZGOt+YrIxBOBBMbV3lqvj7SAgBsG
hwToIhuAkSSVktu/YSm8f4Crg3KM8zQb05XD5z+OMoC0ug/77ElCB+OOBzwf9AhAvqMRTg3L8e9E
vUXWvGVSyT1yMa2yq/AGoIRzU271KxE61kcFd2FRmf2mhaJb7Tn+Qbf2IgOJa1y2QRglNH4nBPN9
DgHZ0mvQj/St0HOWx8ZzFoapVqcATM/MxEdHQNaoL7KQSYG9aRrtOInmHIIcLXvQf+URc6i4CpX+
DMf7zKPVoplX6SlcAeajeXR0eZ3tOc3sO3GvBz6DUglKnSUW8KhBriTdYO5IPfron4JgPYr4/MnP
FmtXs8angZBVwqG0S7McaiBhzFwVmdv6Ki7FE5CrdOQICyb+tTwgmx4Lxz3IXARsbsHXBPsy/uwp
vaRjywSX+YogwHMXW7QVlmOUJf5DNcT0o5azov47/iudWjjITWx08YdUJfag1E984wwQQSBSiX5V
6WxcivyHVVDX1n53OPR1+C5mUrUZ9pu6RTdvP9btzy1+KKvxgqZ70gP80jfi/n8Hh5JlwgGkAIej
YPosSZNNlosgEYAPIHAgYYTTY6wB66Pmzd7cSdgy1wGl6CHn1FqQuQAKVddvnPuBRtiWJIrHLiTT
YQLygEo4i42P/CrUXZhhc6U2cT7tbi6wD/IlHG4+a78v3bNu24cmSrh0OArILpGZcxlbWo9fkaOQ
GaIYFo+rUN6NgUUASK41mlCbGzDiEF+9dRHmjkpSre3cH5Far6a7zOW2spOQTOCfUTyY+9Xd1zei
/XNu5B4bB+L18aDo8XWQ+uZ3OcrNc/yEl+8dexta4yCIlNgL6+ERBqzaoD5BMWK4jZnZD9GmPDz0
2SjjZTnV3jObNi0LSB6GM4fj0+Oti5VHNvjGiF9dvohkueu4O3fOn1+vj9Ap0suDKOlcdXbYfjj2
eKDlaDSNYywQ0H5vHWFLDjpSEFCfYzGHrZ0w6lG7zyhlWCCn6rUw/MPatLgZphtu+swSI2e9dFHH
luM9zIOVobsFrbc2Zky8rfeA97dpYyB1HENKDBZRcFTx5lCpP/ePQQ04//xtu4y0VQ31gHOF+BoP
Qozkg8s8n3llkP02o4RZQ0ley7kFvBYGeo69Otk0IWPQnQMzYFjPZ3Jtvhd+IdAfQs9F8t4nnnMt
D4MSRnTJbHKYlAhfvPxf7EpPbxy7Z8AgBpQEKfYPptcPHt2Z1tv/CMiDHcjpXCWrIk/hoKqun59D
wkcryLrT4dt6Rz3pbBaSZYNGnGngL0l+O2l2W+DP7Tc4d0f1+HBVaowLGrGUPnRaZ2k4y+c3H7Ev
naW4DLVJVAlfZTsKATnYvv9PaNeIKkG0Ci2rk3rl+JPXON9/hi6XO+/fX5sFzB4SvON1xK9M4Vw9
+7QCEH9Syj1I9InGllugLBm1aG0abjDPbWc+8UDGO8mHleBItbFVuDLzfVV5LoZywSJXuro5laDj
kSFb2HPqh0UlZ1vBq0z7cREOpYE=
`protect end_protected
