// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nuF3CGr1kzI4hHXiic7ElhPk98KIuHvtaHhsxGluxzwHngu4CrnlhXR2lr0Z5CT9OO7N7HnhdFJC
RVCeJ5rYxhd5dH9MGpUrWX1zRG7a5YpHH37Cu2zZdEkvdzHJgd3mUpLKisviI8ItPkDkDAEn4kWi
r+3KHFaVmGoA9fRRhOVeAFuKni6618Z8aaNozXrV55kccQfMK3ALElVg7dkos9EKnSpcbiP0TaW5
yndmGJ9uP/F6YA4FrHO2dgyCKv8mjU2VB9PZS7L750S4BlCXqH1ch1Cf5VgkeMDT3jWvnVPo2Vpx
K79BLjTIWA0udn/KFAspjXUGz/qwR2vsw5SCMA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
UhMjCK3d31+GJm2OHdtS+wJKrhoX/+xcm2XBCuoWBDvda6pL2rdMDTGPp8lAW3igQWDt8lUnzEZk
exGCMYfKarEny4Emg2tyfD1jU6PcJg9MsdDXRwzW1+OUFPf+fFX9vrH9tgqADpz2hSyNHE2qkNwf
HcpKx8r3xYInwNKl6LXmOGJXu082JeJwFMsUZ052wlM42KKZ4BWuxPw/XOA08TXon/VOvjwyOzPc
2AugYeiWzNRmz8D0RXyAV3JQl1UQkpal7YR3V7tKu01oUCQAWOVQDDqe+rfFoGJ/hAFsphTUVj/m
85qiaZyd9gjMgREAxeiiEnBHKzjDOZwp4+CHlamPfM/BiU4LtbkIQwRtvCaPmmVTsFz9YaYRKYGu
JU6491mjhXw0Q1QByHlCDTk1VLX4ku9DYWm5uirxhcHyc43T7qSWNBB2tEAEyZbsz+4exgk0aYof
papfwl6+X6TqpYDR8Z52+ukSCTkEunHB9HSs+wipYyl2Ty4pPM/cSYdFc3mXQX9eJicGB5R8lNkq
f3TWlh9Og9iREhLGQ8atmQYyuywX5ZrHo4V4DMOg4KF5kCDFKUofnOXuEbHRxriII8QTIEGthEf3
6rQYm5qqJL18pMPqF4y5b1o1yUs3snC2JsDHVT/Pw6TbIMeHeolTQGMu1T5iKV+sDTpJ8VHSRutY
9QyTcSP91TVsGK9cSjc6ExYUpGXJSJhcWdsovd/0FDwWDeJmK+N2tsQLebHr5Ax/ELU80wSUW/45
PMixsHKUSj6AsEk5tkxJG+ZDcBvqkHlvzVPl4I+eut8+md8piRNQn/lRKC6WX2ef9tVM9MRLOUkv
FLSM6br9dztXjAlM0M60No/i17UBOePP8Nnyjj9w4In5CrYHKOEdD5Yn5J3NYD7oMCWyF1WheSKo
7mVYR77kKvSMJddQYtjcPjcAQGPH+Dm8LWFjPypceiW9w9Lh48l/Ov+VRF8I6FhW+U050RPVfp4+
rHaJo3aCv7jzcrGw4ymEA44SWEQYoTfdTgH4R5XL8KOo4iJsb8wQf/l0FaTHVv0p9HQUdeamZSs7
PZM2XuLjuPsAqV5CLq449NO2qQkLO9jTnW0wyAE8IFICdlMzy01M3m/aWJLEDgAqQns74+inD62H
h75R4skkQVz9j+7b1j34jernUmLTWK4dGCIu1TfnvQkmbS0ZsumdDdrsmwWZnWQgsKOVmwKnEvNP
622WM/nrb8GMKoJtwKciEwD0034K0CpYEXIeieBstmii8pSnff+qCs/VW6TAL9Ahp2rC400RSM03
2A05V18oU7kXFunqzFhyam1zESWC2lKva8YR6vIH3b6ci88cYyLM9zlFoe/Hnr9XLhWNnc/wqGk5
s4HBeFfJKnTQOCx8mDQlTASKYOWCGLYwVGyx5sOI+bCIz+f3R0wV/K9HunFGnDOLHqu+hKwRu/YP
r3aLBl/5I0P33YOy8P7jxb+SdCskt7VmWZEtNehnvZ1/VwmP46dUNTSFtlN/d3alik7j7o71Dt8B
cxtF1I/B4Cy+G7yDKZqMBlqEdZ1Fo6L+wcLc59LkYuqATFcsZoGMwqnyWfBIytotJjJ2DxW/tfYB
Cww7fDUeVtiYI6WP1k1xBI5fpAydTe+L5tab5XNCr31XLHddtj6HczRZoJGVKglYkx5rCcZqaajz
Rs2WUhnwv26jFZnrhDjf2DJXJvqQR2f4p9NhZ1ciHAsMza6t3pcN9iBaVDT31lfF4gLz7gA6NXVo
VRa8EAMHKfeMNHtSAw/G+t2GHBHkbJjTLtMnh6fxRfnqF8sgB5yqZMY39jO59mNqf2abMa95itlC
06OoB5N7KaL4wSHzCXAgpxTIJIaekba6Em7/rV+0gyo/tT18oKaZ6ZlmNPCiVN5Vd7GOMKgkCtHz
JppRqj+3L1gaMtd9R1h6MmvbwQZs9onG5ZOCXYBxlypsKgTz5gNf47K/OP9R4856/QwEgrTaho0M
bk+UmGXSMKGzc0mQOJhO3Gg2Z6CI326QqGULyFpsriqcUUKLdTSCZk5v5BXjlDLY8rGKl6R0yM0Q
7uTdFYs+khpmMUFH9EM4R4AV+MzXlyChH3ZhTyjhb/isfrQrhjILCFb47nGcX8ij7v6+XXbmZAF/
aFXndRtv834iOBWZKAzkYuAABAt6EXeVandDpKjwfkJ7MCNnOcKLyg9+sqoMktE6QcByUA7ZXKBg
fwT5qt5XRqndM+INH6c7OKpUdaFCjfeqpDc4sbQwgOQVZQ0+AFRAEweb2XfQaK5nW9XVwxCYpH3l
tzB8BHo7R/PpS9RwU2behrLiVNYjoYMEuLc3Mdoe/JdYHZAx0rJ8R45pN2um5/679lODctTXG7hv
yYikl7KSfXY4dQMvRCKIwuHpjyLVPIyGSAkSFBZLvl3V+P0Zc3BBtPWSOzOGtU2z9kCPVjS8fw2U
O00PaNSQeOhFl/iZ5ofgnvaL0QQzsXbB36grkjRaH12QCs99YUxz1mQu4/zKN2NjYWgGRM49IC57
jYkkUe1vQZ4iRKsXNuDbR/GtL2Qq7BDS5PqVFLr6KYgWNp4hOi6Y46+Q2kIMUXYoS7O1RewmCPBJ
Jk4FDPB0Fe2aJtufftJA3i/Bh1ixcLzMuBVTOT9kuFlIURy1tPjWZzmJguf9AkfpJrnqeBJgn5Ul
JioSFOt5nz1927mBDUbarh7lhwsjWgVZNgmU2AM+XCpnaGARB3iBD2XszQvkEK5/QRtQ0U0tGbx1
N3oar2gi1TF+xpkfAWCX0fHKezc3hgLyXUhXrImujCDgADZoETUpqDrHI3KuntE/uO+xJMer0agg
wUurWVaz8XrjXTCsaU8kxIWjcKk3JmLLOeZOppL8Nd3s33zrCR450l3TxEp/fpaukjcdGLuoegFP
fh5MwFKqgBorRgAKxLzeOBImXRgpiUYQhEJCH5VfxGXmV4Al2sMqzcOVQvDQkXWtYDP7n4KkqG7q
pFdJSVQETGDjDlUMHNelV6k+THihvls5IZuUG3ZZquk4DuXXgvFmIAAtawtnH13jSFIPGCENtdCi
yclh77NWxqGKJaKbb0AMUolu+0CPoLLN+rRJV9xJqE6rk4n3G37E7pcTC+BOwLs72tbNqUQ9XSVJ
CVKLjwDdb6LYf84Zk67ysXBVPFg7itCIDpwXgLM99rK/NOygeLpEnC9IcKz3S9fLSeyJA5vuJZjD
k0pN3GETccu8N+OR7fs2+Ipab0DA6SkXcG3KIJBz1GRPWQxozBDnWXuKvHIuqe+2zYuirclLg89D
uKCwypZ+a4o7OOLx4NT0heITh1RVBiPafTpIXWw18z0FbrJqGlnvxgKGZqh7SVe5fyG0RwlRgDYZ
UWE+KLkb4Lsmv+zY077S8DPzbmsGZgXZkBkF5nz+WapjRd5Gwgmbfl3aMr5Jcj2ocLYm+DT4rU/N
jRquvdTYxUBzI37TVS5E6pgwzxBC76nyX9JXiMxYtVXDKc6S+dcECvqAMjRDSrmwRy/+LbDtOXtT
/SiXU0cu9JJjPAy6tzl3sU/fDNELJZ1kEVqnx/WSH9sLVj4SrovfoKIi5JLh7Ul4N+JlDnEhnHJV
rsOdJup/tH89z8d8jU0mx0yd67GcLHH88Vov0cIXCmVz08HMeMxT9ZFBDskv60IBgkfDcgnypi4R
CIhZDVHw+HtGHLBGxNZ36m9tLo6ONf/hUyYU7lVYkwkqkcoECNXYxdhro9AL+Hvil89JrugAZb9V
Mf/1jhZ4vPzCCb3XqF6OPdQKjqk3wXhw/jYRIqHEJ0J4jW3IKVlXRp47UK1/UaayAthp90wsaioS
zwFtngNsheYVI/K8rzywOLZWS5oiscAprvJL0zv2bDsYDXCigot2TrI5W0wkDFW+mrGmg2X7C8HW
Uei9XbkXlB6lFyqQ8rUJT+mUJ9ysid1hkVt1xUCmYEoiRqDl5b+/K8mtHvoOSye5BzRkZTo8u5Dg
dRQgiIsfJJBEbvMkfFfcodKl6z0zLiX8WfdikO5nXEDbLPAIiGJE85I/u9MwUuZFiCciAjfqG0kj
dBeGP0rpNKRLGQCkViXvr1ROkn0TuF6GpwlqL4t3LR6Jxho+kno2WOgetGA4fQDnegMRd+JA6/H5
D37p8j4wOxpD99PZuXZzO5taIpDjwqjlfEeiqR2UK354l1t36hWCU8ZJIMK/33n4K10TF+/WWgUF
L5kbrVgN2q9ndwUI0EBD/C+5iciM4E1sWOxO6f4WZQT91vZ4GgS+mgx/Nu4b+ua+sF77NMXjWQty
u2nJ4q4o34cshrRWG+ZaTcmurRwEw2BNL44QwvBAq0TL0J87WZGSsSXA2nhUmHUjbILH9SU47Qzu
JrE3/wYTZo5o2ksfTwMAXq0SA1KQNgiLwbZEwBWM5969dMLJqE+H51EAcIM0eRRM2X2bYhN8FOvN
kW240KwAqFGx2abp3yRP5aZzuPX0KAD1wYzbnvLJN718pQ5sxS5zCMIdXnbngzANDg3TE2KJjfLp
nK5D1epjmvX80GdXrhRiMOS5iYu0SlHlDKdD/lmbDhPhlfh5jACk9M96T1sL+wx4vITh1tM6fXNk
5/XrOAueMutbMtql8a8W5WBDyEix0n7na6S4fkLymnnBsDTaYL/egKECJq/CQfIMF3xZ13GEf18d
1emmZEd1LJzCW4Q7L+JMUgMSuXMXifRQksx0SPI6r9iSoe3IbvJ2p0oLvCDO+HSpTwlXV8LM8QEb
2iIkJhgWLvHBmElQCgHffRDK8VLZBC0xRUU9JqnqA2II8SmRdLxvN6SAph3wKOWL2bUaw7Zw9rK+
hF/LpbqAo0e8xeF00DEd3lMcVEtq+lM47tmFmL4FziGqUkhSy2J1ainExSET7Dj6/lEpIIMCsL2D
rgVWze1U3S+g0cA3z6LyZFckDkzfIacvgOaE6nkSRjglFLvbPTFUqeEXzBSs10h1MkfM/szBzt1B
cTA7g43uLZLNcVybPDVRAApHbBk4SwfB8NF5V5WW4HmA850NgTVevQeZ/X67mHK0zkye3XTpu2wl
YCKLIjLSvHYPAFkDfKluIQ69olU13Yfo1bPlapUQBVUj7gVQtNY2U6JBclKaa19CjyJFlHrdCRht
6PmQsINS0rpIpyZ2XnFKRtF7XlVFky6rvC9pWYQ7zENxB+Kjn4Vx8cHrgPrqlU7cS0WVpIcES3Sv
BnENCIwlFn0DNTudwTGnq3iauHnIvFtHmO4P+lHxYAMelnaRGuf0cseUgkYt4i9G4DoxK69Iq/Sq
1O72uj8Kae7yO5QinSPKJV+sacgs5vx2/X6Q2Kl6byvcSQQPe/j8zf1zQPbP41GscOfgic6aKnNo
6LlRM017Vo9FDLWlYBTztBTcEU6L163eXSdhMI5dn1itfBH9OjEVtpOrLMa8jpRD6qb/SKHDqXEE
xlxUooStosfrpfQffOOgqqhb1ODx696cddXAz44vQATHl/gyaefunJ2CSX6TC7VqW0V5Dlw2JplI
JiY7lFotdvge4pMCTNIgxyJowAKUd8U/HRzt2cJrGKo8n9JOGyLgaeqDYnf/KuEEPfXNR6i4h2qN
e3G3ojoZ6zSVrxoNgnff3fHsTn5qgcR9I2JvQTrdV6f00s+Qg13Kd4BE1yuYDjxc/WKJwbAj14at
RhQ3ucKDPbVxhBXCGeXtZBTKbMIZ1BEegT6gGaH9pUPoLxQ1WW83Edr/kntSOmoS6o5sXVcYyWPV
tsF5m1wAhtKrJpV9uXjn29o2lIz8ggL7lPIAD3U7radwQbBQ5WRKKdcL5nTYSdyDbOtej4jyc3TJ
4rNXfspnLdR5OP+grOfvysCmgMx5yJu+eYl152L5C97fLKewINnc5h4Baeso8gzesXyGwUkF+XQS
/a4ODSujAbQElO6aeShdhRddQyEdUyZQ0px1nZK0Lerrd/kEVI2zwnK/4XvnxVBa6LvZOZ2jaAVs
tjLGSWwAnJp5b6LaE1zVIPkX87nUWZRNVTsh3X14AAkq5rPQMAq8OMEhxlZVPVWLUnorIPtuLQKf
5F2zasepaDMlgmiSkVtCARQeUReg2iLq5JNLvbty/iELZUIkpyQgJXyZxpuVch0rLyxj7f9JD5Rk
QHKCfpkP0/4V9xgy+yuKAckvMAnq4q+j7O7Pxj48R5vdcwzit4xxNNnR+nvMgFGDyvSKiZLP1D2B
235vGs36JQC51nBEX+GeT2jF/gPATNazVY81u7rGWkIrAM17E5HD67XlpSWMEJEsE1jL/o/bKkF8
3KObC8OTZ8WhjFoeVQeoyrFQnsXtav83Sar9QN0hoyBPCmjza+E/FQDJ05+RoPc/rKUHxo+i5kzf
Vu6SB4YhAFuQ6mVTjw73RTf3F45qDyDhRr0u0q9nylJOFDL/ZuHpwgZr4VaA6LPWOQTebhWJAOIc
oUOD7wenav+zbRAP6r/0xPyRxChLLKUH4hXWbaxa1F21Zrj6Xo/X7tENhlv6KfMKt4KnBZkgd5hr
UMgxePP/Flqifd94qkFhpWamdfXN14Nb0nT/PoEG+PUPTUbR8wKhh8Ax/XL8pp2JDmG1LEK+lKMq
4VQq7Dm0m8B/aX8WtZis+OdY63P/lYPUbUISOCixYsG3449xCHQYEPfFL95bVvDcAtpLkZubjVnt
KjR8BXzp+oP0lWdceX9lNRQht42Hj6fnUeH5dV5uv2mUyhHsLPHyd33FCfRXO7KxoZDdbs6xRRVI
G/Nm4bwURbi2wgysJk0+OKhnFXaPJtmnHRinZ5UG4tSXHHPyImCFVAmvoJG7sW/NKKzv6mZY83bL
ntvBr1cOiV/uR5M6tvvjSfFSy+uMNYwixGZm7sJCA29KYYhcZ90RGyWB1vU90yBArUOB4P0N0PAz
IaeOuTbjEQ7a+4hZ6XY+oTHFF8eHaTfoZTYsgb9NDLnPSqESpkGwBdUiA1DAOTgrQtU0fsrLUxuK
DPpkYQqwK790dAuf9GAKWpBeBFM0meS6TcIHSYgygIvumY5b9ZHPeQY0L+hQ7GgLZP2O+mkWoQUV
+VMhFPbn/KpU2OiRR/cs3xgtmQdROLAW+iMQnf6tVhU8X/EVbkSDSZzMbHsZ+JRJqBFuVM7Y0JId
KlvkajUSv6Yo7RkenofI4VAb/EZ3hXFpKpKgsVFtCnUr9F2f0d6f2OeV1KQkercJII+uTam64SX1
i0cDyVOTKrKVwIcvFs9BTGCBOcz3wIagKzRGIDcL39PMU4D/RJCVAuyYSV2OUu+mtx8adGAciNAg
rif+cExvm5myQKUttQb1I7m6G0Gr4uCvhHi3OidNaOTzZbtfuJ1oz+XbB1dvEUoRNFc9KgeDFxHs
sQRQ872A2zQqWM0bk2r4wlvPL79l6mw69+rQdsUIHRSBUQa4z3AsXxrSzIXpsHFIAhKutkaxiWEV
wUaBydsh5dAMc7QBPaupk5Kk2ImDNbTuYoMsg/6E9PeLcFciZsZwjXnNqnzE+ZhDdGQm1+GRPhQm
nAwX599EkoTuRwIBhs2ZjILdXBlVfzGneql7jmfdPMXjdNvAl/LNvZX3ZqF6C/w1YTyXWhM7l28k
V0NCv8d4fDtbE0vp+m5YKNr5+GZeZNkDjkc/yE3OpP5zBFySu08lQGHXaYU8vaJ3iAcdsvpgCL/X
s/70UzoysyE654nCN3RAG1QQk5FcWbVwmQMkmvkhT4Xd1sPCwkCl7SIFQCzOLjZHoyl7HvcLgAsd
sqdHaBi6B8HBjaegy4DXSCHKCcwb6WFjtNLGL08OHAtPl/M+QdzdAkgVLuR3ghe4yLdOWH1SeZVg
cbK4x+aVaIZqkfZEiEDuoecvPyzAfPjRNv1ji2i6ytqQg3EqW8grZdsSxeUl+NwQL1o3ZQcH3wLa
Zg0kj1E7O6MrNvEY7qxrK0FMhiVI3Gf1vZujXrfpr5CGctPrxzXUmLYcBrbc+Wdgdh10p7KThZ/D
VZVOUNtwczYOY5yVOcN/aNbtpR22niIN4oRtAEJvigUjjd9X+6bCRsEzYYlJeER9D59w3OcOwpR9
EyFzZA0TH2BMdgAvL8cuSCWBfMPUTCntbV1quk9n43JULpzjZRA47egyAWqUlJ34LeL+2R5a0i2v
97HxMTYlHaQcdS2ruA7GGldbfaOeXvxs+nPTJphWYelgHPRmahC70cVMZvLpl74lUksxbh+BOCg0
ZrRb+pOxNxcdCRI3d2z1iE27Jh38SLDfyGM+iBiPujwYDD8OzAmaws4LnUfoJp8ft+wsSWd90pma
IcAOldA6f2YDJN95ZH8UtQ8ePKlq+oYA0SfwR1bi8NLOx5s0fRy8wMxHnar2m9RQrPjGXhaT+Xy3
uliKnUNpEeJzRP0ITWNEJulf6RwNkkeKowS5VV/MS+d3zjHPj9k/Au6tbyZWkcl56twR6SXOIcoO
8kDldKXNUFjN7mPMR4cOrn0KoEj2WXiyRv9iIUv770nhPlytwpEk7rh8GamGoDLJiiC24f40gDlm
8MfqBIT3v1ZrEd7G9BzBurKj5BnWHFOBLM72Cf3HffgO8fiv/ui0GkqRx7TD9MKnBuSt6ebeuEmT
ZgYE3mA1/IS5DVlVwq2YIha02L57IKg81gcnQuR9B9y2OE6vcvTYyrlxGI5rUj+V3UvEWtZ5oCL0
K1ChtZBf3yQCKSXV1zDhQHVvyu9LB3WUf5g+cDmXydM7YYha0/cYLOFvRKp2zlIo0DzCEglPlJZW
94yW3l3HKBOcaochTpOHr89DZIeip7K5VdTjzji6qy2Dr+T0GEXLsF0RVfW7lM8hiW74B6MkLUpX
1oCJi5/awNEbB7gB71KNbayCYNlBxn4iaAtrFCGqkQElgOX5XfXKUp/17ETMGzk54B4lkhJ6MkUn
DauTJ7R4/Mxw9s8yMayePIHp30HqOw2flODJRQZ+5c+9kjetKhuUoaMNz1cjwu+0GIkTqNgzGWw3
g1zI2S4GsJhnNeyXa/CHtBCyJw16W5yoXfc83obZ/4Xo+14N8esUwgz5qDR5mdoSecyP4FY+bRb4
U8VAKmYno1do7PWSLTSrq3XeRhyBlnHqg0+8DLLoa/8QoCm5Z344/rAGhSQlFK2XkrRZNUBWCTY7
uymE2coKWOntKkmYD2tKNTqYiQ+c8e+dPA5/yFrZLJ6pYfr2J61HRj58vQhDkcAPlxE7GcA+gXYL
43ASjZh882/lqPj7FFR0ICeVielqYB1cHxO/hGsud2/oW4vsGfqnDUOZnuEEK8zVzCQE0i3G0MGb
aXFzCTTWPVwGMhnUSM6R+MyVrKcdaG8bmhlWyNd58ULQETrRkyrgIjRPVW4ILU7x4iTEeg8oKOi+
lH/AuVwe1tpunj4928fl4YpeyWxPuzVWx3x/Z5Jc1Pva7oRQVNirm8ZoMFT5v9nvp3y6RDG9IStR
jPH6V6ec261TfhQjAyO9v53V3arGmIAJRPiwTdPhUHInfE0Fu7sY7UROUszYsZwBi+UnqLnpMeTu
0FXILZFu7icdE30Ur9t++MeTHep0VI3683JgvbaiOl6V+vDDnt5kozJZcsULWdM0bqVzcCMvxwRN
cmwknpCX4kn+rZC8UnAoT13h7TVoa6BwmWvwiQgQviVz8ssmJ/xGmDf0CHTY9Ji78KxSvs8iT9ol
RGPEUjOTvbbaFwL3YpXdYipa9tlZH3WdPCcSxKDde42MrolfX0713GHVC8LPEGnVt60hf1fAHGg3
CMAPsjKm4McL2+Gyyb/4BteKbA2/Pf7jplcdaAY/aRMDI97gY2knOBd1sa+k0hQ1Z0AL9l0AE7nX
OyfZrm/N4Vz4Y84+s0uLwuY+QjgT+0AmMEpB4GCGqbXYF2YZuqkLmohRVX6gosEqAshv5jQbep+A
P/YJa09zXKcCiw/bEdez3kWdHfN5kcIUKJGykhk7eaxKh71W8mcmoBUG59bxfWaHjZ71jSGJ/7tu
9uEGFsBBfnkhIvq9ZafWyO6uKL/ZZ69dzS9OO0b3TJKpIkbhtlmHfIJh6P9q1DSVJllOUD7f5mLv
zG6BfEGKLTmhXlGexw7fih2CZe6lO/4tg4YUGTxZ0/4QVSDjC8TckxuYH699XQbJffxNEilbi0x9
9XhyfxK3U1zq68+RA+v7wjRmqDNF5rNWj85LMNTh+Wwc7Xc/4iVPxph8puAXJi8xGYJlV3BqZS2V
6slxe7Or/w5+M8uM24UkII26MVLJpNa3/blFrMeRkDYxENQPpyNouJSymKK3WXLPNAVelmlQNyv/
olcwDiUHC5aTD9c4OeaHENSF6Pz14Y9a5BP8IL0JFEFF8fRPMYpJA4bMDwdRBKFJrQ2v3Zp+v9zY
2tmE8Gx0266Qt/N/ufvC0rY5PzCTE/AIcuj0HoYGqtkjumyKTfbXU6vv9gwfXgivpT/+H9pd2LCE
76yovSwMX+zxdF/W1Gg2PCHuizaEqiRpFbxGarNQ1hCvf+HqrTvYRFEcnMvlVSqNwwvbj7nxkxDj
xjhz3+zK3g508QXms3tX79iGHOoSeyxkjHDLH6B9F0ARg3ACPfCyCAQrkY4S7O+PK4NzJCCNYybh
/MjrUx/IS1QI5hkUxLKBO+I8XPfYHYoMUlXa7gA86ESAJsbJ0qmM1kosdNZGKoXWufyvPcjQh8Zs
/aEqIiCtm6MNR0QggB/oNl9qUFHufk+gdFEKqsop/i6c55PFRMXwnnC92PsPbmmI5lnn3030bFbb
P4obgy9PX63alZfdHIc+PPyvuLnAVBonctFwnUZLHGiAwLovbeDYR1ZGGg+Mi+QYMPKX9oMBlSOE
panp8IkluSQMTwNNeiKU7IDYg/O1cMIC/a8FWr5RVeBx0VPzAZa7M72iRawiTBn/UgVU4DI2I/g3
kJXrAqRvManiu/yNsBkHJCB/nplO8HWJN0TiKqVs9Ch3PzXB2pVchYZfVbfAIkp+j/iqaDbaWQGD
J9ctGA6izSODpJLTa3HNX236xyZtv+j9gy2QAPoYQS0JQCA5MfKi1q5lNeY9sJb1QpMdmhoKE753
HqdGhuN56ErSLLbko2THnXGaiTxd/E7H2YFDaBe+uAkrAZYM0UsgZ6PTWmEeYKHWtMua8KENvLjl
0bq4bm3xPDU/hwpxBkqDiPb+XuKlf1y2Jheuf2L7iZEBP9sxC8uBBLVzal6PpTOJHXI/37dZvuYT
wBQSj7b4bg8BW+uo2krut3SE5tzkq+HMUzpUvybglyprO1/QCiryKOjEFbYxK5ivKLARVLQSzCPd
yfIHwet8Yonj/9M7Lu4PKUd9Lx6Mxn+6f/8qC+Uq6ebFpXdA7tg953yGnfWgZ3l1MfgyW/MGlxao
2K9w8SLetqu86fonSCOYeQrQQ6Sb5DRGXOOlDMets6w3C/ku13Fd/cUSnqT9y+l5wwQ8H69BpnVz
7NsOhV3VxirlY16ExykaLXaFOfBtADmtTvWw/jBKhuzdIPCrXoSUwjgc57hdBe9fSUr/SJw4c//n
bSV1gFqxk+dUObjkWEFCOqH2NwxJD1qVJWbRneRf5AgcgJ2hyna4l10okpI57RO79CecVItADz4K
YvTw8VG/gxwAjmt0akD4vMEYJGkyMBtbsALi/mRpBXAm+aTdzjlRGW4trGjDJbyTx8TkYe8qIIVi
vlOXxDqMqrdln1+fUdKLTzCeV92fayvdvc1tt3yw4puJIAUDBG9VDqyHppRlfVMVLwgvG9SIUsJy
RmR8v3gcTzyKFygRxO1pejoDgpY4AUtzAuxtj+3HTXUhtUaiKI8CNAVFJa8mv10v2wp603bLjyoP
p8RPJkXZLFLNKI+VvbmL52mTSJPOdUH8wVtfAgkcqbZ+sIpcttweDgZl+kj2wkk/JxSxU4yTKNq6
DjmQx/YiSpt/oAIwmEdfztiMv5OHyiElRbcFlFY+sqonn8wLAQReTNrzRWeBA2eJjHU+uq2IRd5w
Np18PCztVuggBM2XCSDGte6V5Mh6hRLRQinENYtJyIx/cFoiFzPqUHs7m0ZMr6gpzNIIFEUV1t/0
W0/5hr5laxVmBRX7ZU3aLYLHv5tJBC+0BQcoQX+P0ak3xDrEu8AP1fOZ7uCC+CHKmj+u87C0G6wG
KCDK/JuqP5JVfXwm2IfIDpiNbbPr2jvT4QqaemXBnSCpoIO/CSqfPztnxY+3x/0BHLbS3Qyd5yHv
3EhHtXGAWVRwbG0FwIOTIbhBk33VOqmfWyqBT2TWvUGJaagBb7hcxevXek91Hy8P7Sfo5dXdVmih
Ii7Nb0gmqJ6y4Jk0Lv8q5o5T2HnjOuh0eYft2ePrhkQjxRcPi6ETuOTvzzlElj+8md8igWtMW6aU
P+DhYCF00esYTXs15R1EMWh2QLvCNIqdMv4EXB8AstntFlbjXipd/pAFlU21XCfV21gWvIGFOwX+
r7ewdwswzEndJXVfaUUb/JTvMK88cLQYBf4iMFeoQPGQWLQhSuB5zxJiRe+V6VgyM9pCMEbDayST
OtMkxrnB/OTZSMXsj0t1bSI9nc+8Bf6fbhkcYdWIJBuFAXp2MK/X0s5PPcYumbD0T48XVFw+8l7y
oY7zhx3YBsFRUFUeSbuh+Iaq2k5uqmDokDSu42oO8HlHRQAlgkm5kCx+ndszavZA1346PWtiPas7
q1skH8gr1+7QbnW2+/52UYg7aLIw5UodCXQ8fQH82Pog+jC/vAwGHRNp5Qr0nQXc57qZ1d8ixvK5
PVwyNzbbdfghTRnv4EhAB6WPgXEvHm3gVwRRDOZm/VR8qZhA6ULOT+UnZe8Nha6Ud++I84vZsPXc
tYG5KCrbS6IzVOceUtsdCItnaBhtuhIaQlA/8JojgpcTZYt2UDvuWsg8SBhO1/F7EaZeXh13YUNt
IYYYxhQvVtCPB5UfA23QQjZTtxasQCDt6AsBqjk4JnaGB5IUwoKcaeeY7rfuTIaFu1Nbpdmxx4lB
3P+8RkyVb6IR7xciGDAYdLm5wyahNpVNmh6kvjMba5QxIJrLOGhgfdrVoNGrAKiBqUZujBZmcA60
KMOvMKxYFKrahSCv5UvktYXlFWFMaCn2ifFjp8POUlWY3evqKAJG7N+21GeifPD27OfKPW1y5xhb
r9/3Uk0vORKfJkozRIJVLahAmr/lZBNJLv214e8KaUTEYVFuMyjx1ZvIaO1onx4oEgf2vUXY50uE
BrpfJop0FWw6ZWHrlaxSMjZCPk+d1KE6vqJx9QGCbDZrfgnPMWc2mZ00Z1iwW+DEkR425W7cZMrF
TUcdjN/WmHrLvzz2udZlBu66mDKEn3bwv2bXrrEHs7bexASZCW6lu/eIsVA4vBDGlLi1V9ruv6Ti
9j3Vo40G9vda+FdKo3204bua/fx+kFTrYU12DN7SvDR9ec2XqZfkJacodu7D1niuc+dvHa8K/0wB
elkGMWUnKH8dDn+EPvL7nIcyqhNNG6/6n2+1SZGprWi41XRaloA+32As6c+ImsmzfxYmnS9G14jW
taiSGhEBI7Targ+hkfMZxAgEI2xrVsfpToHAZztUQQ4tZgV4Xx/gvnG8chW2V1EuCQAoPjxJugTt
xI0RE2SS2bc7QisrRjj5Bb6yDiB21d9qz1g1cTWPuKtlr6Hq8lrcJ4ddbGUoGffg37kU+98A8q6H
xbc8rnY7t+cOxC0ceT5hUQMvdElCRVUEVD+13fJpbH/ixeUhpjIdDZR90M7NOGfSc0ARO/HxlR+o
KxNJZJftMI06O4MqszWcqhsISPjxbuIhoLmIvpdTjgK8Mmb9eq5d6VzlJXtCy2yKRLaXf0+dg9fg
4WSRo59E3SP4uHzSOLUbUAna6yOgQyFtFgBiB7dxgd67vvqF9SCwGdrY9Bxqs9/9++XA3S0ORykB
kTpjvB6IvMFok/wr++Zjb4HzzaYMpNHQjanSj+VtRBk7NJr2PwhcObS2KChKrubIX7r5XkcUyrYs
fyuTjH4DcmErDDS30LVdZBhi6p/vVSHM9t56AekM5AIJ1yjIiHsgbBnnCZ2ff/qJhfsEevb9cor0
1ULb6Viuf0aJR8uGxfDoZd9K7SbJuCfUrR3KtuVNyfSq/7r9C2t7Kq2FrZeEYvgVWI069skYj7Io
a0Ktf1juJ8y1PzNkpmVdtNua7lOVVdKEvbNuFw8XOY5AKFFprpcXdRx7y6/1wnYgJptqEZz6NkMv
bRUQEUIFX4r6V1RqyvL5xvncm5m/bAr6kT+asTkXnRDGqeBj9KXFy3iMFaxcREzJOaRX0DtyMWv+
cNep7QaKHmwuLJmmmHVaNVKeTrvaw8s4x9mzyKte8cqWwuIuHqYr9H5bB3sMdVVQQV4iuQSJDq+n
vgkJ+MiD0CwWhJ7H0h5QE+v+Ywc6puOyDrgrwU0vglAjK1P8Qp05cXzbEJsuYLiSKBKaudnJV0Wy
5JPTm6DJpk7WocwDyKypTOVmSmyPPfaw9rgwmuJEkUC8K0GCYR6HzRdosexuFdL51pMwQIi6zBXZ
YAbIYYZu4kZMINX1JSk4sPtbLaKfHl1/Y209gQ504seNZlAKCnk9QNt6pnqWX2Tm+vilulo/miWn
eqaSAxuyHnbM3QTL/aiVlD0402F/I6DnSOlPT6MwzvD+EjdKk6WpB76hSLQLhBsueRuu8jlvPdZ2
7UJ5o+W0nPgUXnODnqY+kZsikFZ+LXSc5yhsphxeOZhKEd+sA8nMA2lXeh5bk9VNVfs70Mo9kD7K
ulmhG74GWQkf39RF0jYW04eLC6J4fg6cK9jzXb9du7NAfTB3WbxrigHFEFlVTAahAJiwkxR6Tt4y
+ZOxBs2eH5wb+gWSLTuegGmjSxxyB0sw3S3/2jdyvGZ2UO+TYs4KwGVVZKVUQ1VsRl0VWaH9hUkf
L0hdUwF6/9YygPChPttnma0WstFCBd/ccP6Qg16MnrSzbaO/HUOBJXke6ZcRoxCvIem7kHMAcsI9
xijwN5QqXVN8Z943S9s3yc0BGD6PN+ZyNnuMi4SXOFbRy5nLbMMttGsSPVwejacUFaNQ9LTZtrip
tZST5tpQxdMLktVWHstihVEmw0HFex50dJdDr0LMHm84EZXLVg2dfCeDN3Rc8QMkX/WK2L09LzkZ
zkD9njrfsHedWVMpn1O1y+tWGNJCTZBHkSuNTC0jJjnXSLkTH77Kk+iIkPsWdRNFy4LWJFEyYCm0
QpDfQ7gpJ0TSqadoMr91H61+hpHqMjtSerU4z4VshzBR+EpGJlt4FGaTWQkLKnYrON8yD+qDtAQE
P4MVZGz7b2tCXY7i2CxMWc8C8aJ+yfH5hdEunVmu0iXiD6hh6ic42wl/G3i5GIPrBcjYtuDKw2b+
+y/1/s7HO9L11tklVPsfgi+P6ixSpGCv6gmJVHIQV0qTmE6BoYhIh/JXVdHmcHyEAWCTT2719jpF
jV1465QgMq9Gar1VfeZEt0VIPbLkFtzyQsi3b5iGAZHdAUq395j/it8VxtbhJG2IZyMIy2fopPZe
+4aDNzx35e7b+5yCzqiM0oAXjxM1jQDhhYX2YYPMvTWbBbwoqne6d/PNxKDq6l7QCTx+EqGOVVH+
DxEmVFyzHc/i2g9NbIxTTP/g66DHAmh9T3H5SgXq2zPQf2+d+WPQBofYn8W2PFJgbbhbkVtpIM+2
X+qm3MSvgkUrUdqhebZOHIh3Sx3AH35REDfNytZSIw21IMpCjyMtp2w4KQ4UFpMSCz72+lJuI5GU
6zEiC2i7HfY+sQ+IWKGFzteeyEd+P56djvddksFCiFPIiCUqbAZta6I5z1KPOWG/uW5W3Vwvgdc6
ynVaRoVtFrIAYlbDrYyD57FADl0PEYzfsATwBADSFjBKHqWl5HcSvv7eULGWsxaYdYlz4FmfCOtd
fcjlKGNxoQlPwSP82TPcq8mJqr2XLrwdV7Nw9iHDnjd3L3WS+PgRT/dbM29deQYavidmYsqjiScf
+u91yrWMwwB1lk2g2TozLBH/XJGoU7g3hkrvpQ3cEcXckZQ35QeqgHyKv4DT9TbuTDFEAxt1bn/d
M7RO0xrniMP47dXpDDiu50LY60A+2gT9XLyan1wWjt5zOY2kOmYPSTEE//Uv8FIaYOszAJHEMn4z
YSDjxsbpbhAaikF/G7lPkc+BaEL5YQFjfWao+fSZvlALzNBI1q6Xjc+duZKZEAuX0Sar6HCIYNaa
FlobLvwG34ZgAk9ckTtKuMQQfNRjGa53rqc3Vo3QMJ4GDII/Y+Fy0xql5tPXWg2nDMGMzmqom2dw
jvoDRakB93thfkR4YGp+a0Eb1wQXpfSu1gpCc7Hvfu+pXbK1b0CiuRTm3/ZhNhzmP9PdwH8lTKZB
jKmWfhha9sxf/zJW6SZymQS+QvLl2ipRjN0EYAxgtJka6O10bEARvCedhoLv/vNf/obUC5hv1AqJ
dzl8LColGyZg+yGoz+piygYje1wGTfBXojtjCReXpG5cF8iQXjnxZeakjx38oWcbz5dTx1dhdHSI
b64Y2lOp/S8VUPAUkcQWH3cH7WkEXp6Pw/7SOPyoVrJS4PDIQyptdPaB2qD9Kh87QvvU62kvIbIs
jG9GzAVD8GLvEkCcX35nh5hSxaizEeumLzNdWAqFwfR8dwngW1XpbyTScNQgNv2C73FvbSXkYCQs
Eidi3SXdD5XKv4PdTT4dNkXKIeC7IwNZdZFiSsbf5/n4G7KiXwFq+xLsYeZRaBqUVGFFR06W5Ug2
4jxHuvuRmG36Y/5aUgNpMDaEKIwxDciGwk+N+RgDWJckjcJmKxgAPS6gL++Ep0q4IUhQvgZC7qCZ
Ljnh/uYkwGPRBwgrJ2mXpYau7r42FnMZs3FFQLwtEeOptKa8ZTPindFGHrxz1wphBRY5uXJJwhlP
ugWBG45aor3gfR9t6agJfrAzoAPuedvGrFj2Xf0IydUZ2/9weT3nSX1vq4jyxgCDlhmbbAM3fZx2
v3zbp6iU7S4lBzabryER5UQc6GeA9gNep0JwYp8bYkSuaJWMj96LlHzO4M2AlyeObFXDdvTM5Gzr
cU7Z+QefByX9Im1cepWVcZALApNbslWMUVn2v4wpDPm9sJtwxNAKzVJ+iLtU2vLX8TF+LLgg1uI6
xCd5ThPE0t25378AmKJGoCLlr7qLu2A9ns6esWX+dsWCpTko0pu4TWvTO52CmAVVayooI9ligeky
d7FBTAwCP43OcZK5JnUs1vRrZRt/X/utq0zYnsdANCfYXqpRh4TFmAYO7s6lQn5HaDhp91J8tfV3
G/ZcwUxHjyav9i/YtvBrtYK+HZcfU73xNCLFh6uHs5I5Y+k/TqDOA1BJTGN3S51xt8Y8L7Amvf2J
rZJq51SloNrecOFZsR/pw1Gb1fJtcoLVFebqdfbMjafF+HvJINp6sk0j4V4fROYpAokw6Q/DmE+Q
STPZfQaELJ4WfOH4xcPzkwSWoSCeIAVAbF4GZKoS/HtqAwROumSrf7EIBqhDKeilZChLA7SADB9U
qCF5V8xXMolwEcO1sUJ5snajlEmjqRlZstkFYAGg36jkWjKBbwYZD7QSahoT+bZ8W7ujmgH7fORH
i1GloHAxlmmMpgZ/WeEyUgYkyIiR7jxcBSfgoY1CN2q+BS6wCBVNmvRSGuFQyXPIfHlydqOXssHT
lq1MyHa/Gb9u/CGKskoj2VzXcCYHyQ7JFdDnDVnXB4AyrtBMtv4ynC6wS3b0VlC2EZSggfTorvZI
xwPn9fwBNaYZfwG+CiiFZysSOI9/CnJmF6FxmlN7RajqCgA6x3TPMRA+f+osAIFgArR3UcWiI4sP
B9AvNsBoixVl2lVVXNBqGQ4/RPOIrvI+wi3ORiYmehS79fGEm8bGN7D2RngHrmI0g4PmTu2gNmQr
eh7IiEjkoGGisAQ54GhPVloA20DnsYrrFxb2AQxkpn8CXw52Pau8Tocci+IQObPsEtf2h+irmxoe
qnxNy7SJ5x9VuaEcrRdVMDsESv3kXh9/MT/yIHzKkGCjN+2YPUdzwB+4rUKrigYC7Thj7jHgfWIW
vQKIyh1UGdbObNJ91TdnZl1bIJ10LQ7AHWVSJ59CzN9x2EEeSYU2moQLT6of3GqlG8hcKCvtKMec
a7kS5VL2OYrEUH8nQzM4tl8MBfHEuSBhPnh1nzftRBYViSgsE0RMRlnyLYtLVGChcKIxMYGHqOOx
GlIHAVyc9t4ELhb7OrfyjnhOgYTKOScHkdlIb7IvyzhSk/uNdNP2P1FYQ+VOs6qMRi073lnTPpIR
E20PI3gc9KDIjTWFKWAAO/QCzUFovofusc7zpnnEk5MFe/64eEFczuulLNCxfuIS5TnSbk8AMAGW
sZ808eX4eoNprbjPfiASzouxZJmPqUVl86y5ILOLAKA+MLsSP3FvS1JOqipaGZb1wYQC8WT1IHNb
gQR0rvW7lqDHv8a1oL1TvyzYvy8t4q6XYYYFQ7R9v0fgUL9oBBvktq9IUerfWhuMtcLHaFyJ7n+Z
QYbQamEOjklQzYIhziMtJzkPtw6hxsZCfkD/9bApMsiG8SKdTC0RgiqLN+PPt8VyijMvyyrwIPWz
qlpDadvQATOPC7O2KQwaGhhWY/5faizixHmEb0rMhEbAiB8nYAJogaOdoGMskOCRMkuttP4a495i
7YPb8KiePwVQY6Ni8EBN+pUyjYwPvRNq0WednU6G5PdNH+eVMXTa4lPcoGKduEsXLRG4ZIxR+fSy
MLfZBdI74jm4yfex89b8UiJFhioTUMd30tYkWwcpmkrUSsNo/CQNF8CY6B7YI2kNXiyMuDVryYi9
XoMMAns06gEXf1aBt3H4/smnrMJELq4IEdB/hcBMl4vOi/Y=
`pragma protect end_protected
