// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lKbZqNWKdDFU+zYsPFsvzkGWSlik1sO763jtVNz1/HRrRL964OMkuos54xGBPhYy
Duq55cZC19obMquffGvUT9tBmcTpXUMwERgOfrA93j/R3ZJrIDe44nZDf5qLnHwc
bBa+2Vzu5h8/jWoxhPNpw6KC4eK4520nSi6SiapfDSo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
xfRps7F+fZMHiHZc7IrVoqCo11CeJoiYAP0SFs/aZbIWz+g6j7f4oiW+hCOUEnMe
JdTdNGmQidWYeD+iyrhBtvbAbhjRoKpoRmhKuDmKz8M5cKI+aGCGxAauUOsdyTLf
SnVTVmFeBJMpSJbKVhpjs+HR2+BW8E6aGb1elZlMaYBctLbn0vvfpHUKqOnmiegp
iyM9P7A3xB+foGUvIb9oRVjTsvFofwXzxxgpaZXrgOqMNjKE4QV2r0O8Dz0cT7U4
TFTExk0UAlGmFXbgJi6K1wWVfpXZGffzwvR44W7a/esjBWtYxu4C4JQhGZlR1g1S
hGsy51fjufc5NTVci2bMuJvlGKZHTUMKlMmucsg0pGSYFrjDp0XJ1EEeUDuYZ0Pf
lFUOwzkFw2aPjMayD3tFBQkB1Ii8Sd6+7xahA5EfhqFeqbCu5jI1GS62YNOJpC02
SVxqK7P5TfAvZ+h+ZVDrxsL3i0hstQhw2CiV2xYypKu32+w/qIeV0iCahL68fnHP
5sJBLwBxnlVURJ0E8ClJxjtP6ovELfBjqS2lD/iTnmBUhC4tiIMweh8L/POSR8et
Ii7LPtLMprwg90RTcJ7KZxUoToWO/5RzPwrLGYkznlGK/4vmY4Tz0D7fwZr8P7q5
sBNf2mx9Xsixbj2OT2Ujv/BkYIMcggcRD49ss1httkAW5Oc+BIVOMsCj2ii5BeTE
+neKIuPozfc0PgMxDaCIBXX9qXOq7bqhjJpvE1wlURNCElX7n3Kp4vHAAAl2LNnY
qmcahWjasNy+Nqbc05ErVDrCA7TO2VZo+iP06UZB5VCUTvacIIiRVpOEce8rAWAY
hHyrmL2JimlvkAJU/TyG7sKik+ptvX2ApV+9tIyWmzQCwap1i2cc7bT5j72dvb69
MeZx/2CV5hoikNj9BoknbaW+12afQMFHRAzjewVq/9JKGHWKHPp8oADjruduvhLm
iWnlMZLDGOKedb5kTIzVrj4VjJ2bdeOCsQncDOG4gCcAamCuZ4HqUfZV46TB3tHV
v7urcCHNqZse/PVbiGT4eNS1bnUk9CRwpqk06HhZnBOvP332Y3iwmMYiMXBmPhiG
mSDb6bEzZPwYu3b3Uj8g9/iS22i1oJctzYJuddop9PRFG+3ysPQdDeHhziXsGC+Q
s1Dw8+qy7TRCxtUmD79sQkpPlFnCkppOfYqv1GqcLhNKZcmKEZHt1d5/DALWaEiZ
Q7v2SbaPt0B/lGRMf9267bWddeFs0hd6voC7iyqHy7qdwMPsMuQOeJtXbgN5F0S3
hxB8kmt+2daNfIcRQ6zsJ7euTQUou4cFWm8/zIkERaG38VdnLg+TnwlL6QMsfxMy
/ESCV7ssdSznLCWn4ra5W/zypn0KPj1Ib+RLJ5j2tJeRNb5OO7PJGPrr2gr7s6vQ
UP2/zwdqpEPA0bo28sQyKKKJhmyCqu8ocD9FupxjKGWkXN28zc8NWmEeaMJR9kd9
FMaUXlhKVFnZtvotjHc6SL9g5vRjVXKuQQwSIA93psKRy8bavgH9lVrPoi0YHWzq
206NTC5TU87jPdJlRUveACNJ+I/NYw8zL13AZcPMADOR6UP8QTintRJdDXv1pGzI
9fpw93jv0gdL2qSF1vLqpXs0iHXPiHvCr9jflWRo8MiSjAewHiOe/RLYYtpX0nwm
USI9KVnAolmTeBetOvftX2BTiB70PsMFkDn8YUW7ywynXRghp0gJBtIO8uVheqnQ
ZHZydXbSqR0u1tlyerQbVvenMrIhi7VzJX9ZF6EDERUV3vSKyb8k6WpPB0wtVxZ0
frymN/SAupvHcz1UZ6aVmhXjqis1c7cNepGFh5z0vsQHvS3r4erSTlMRwJIYwuwH
0EWo/Nksnx4DDveOBVwQPPE7j9m20Jy9joA4ewEQ/wcyGDaN0g4/3j4xozYP34Wz
SUYyoo2+hOExha4oc8OiVGLUbjIKI+GSVjIAlRfKqDMWHDCN3Qcj8jU4bRAojdal
RWROjh0fPvZsAOkAK2tEm2vYBxIATeSsK/iQO4stlyjhc5taZ/5PmlBLzNtaOv6r
N/LSnfZYo+cPvMGzV3UTAWJZmDBrGDYBi+HvaynwCCft3RH742SQ0A0yLFc4baFR
I1ACN2i1EjkvGIfTbDkk3mUZlfthhsIBLuOapz1ISqQnzLUw2SN5JQEXGXbdmAsI
NgKGWnNBN23+3xGF562J0jLsZlBoEfUbcl2LLtL2lPJMBr3zAhULiexAQHF2Vljm
O5smkdr0R3n+p5hjSWSvdaQdLGP+JH+LhW/XYG7qVNW2hC7VLEhFp5/N8zGE6xjv
WtOlYeKptcOR1dgxsU54sSVNrTeTHScD4TkzFPI6oVpDCAhaufZpxfN2Mrl5lbFA
raORdyWhCyKLCDil4AFq7P+pJw8y6PJTfGmjRRYD3O1hjQdygr+Lsynop5vJzTMr
eZ2FdHUl5S4dNgzY4vc71jwSnsUhjuTfLDg4W2jmI7/mSzVdu4ktcfj6ff768WGc
DK+v3OVI4OD5zZE2pru3Ifro9GwkLPLZGFmPB5e9umoRn6J5d8sxj612gJwG/fzd
ckTv6AMh9j7VFktR9cAh/UD9bOWW0AoA7cMjvrhf2dPuPXeutBsgJjnQbBKEYJj3
U3GwBCr0Sxs0wSDb8F+GP/OoXNP72dXBaq4tyd/rI/Oc73y+haL96ldHZmkNotRY
+WygNTnWa1y8x1QuQiLEdbQbspNfxuzp+dX+EnK1KvXUIIRwxVEhFwr5546oWKoP
`pragma protect end_protected
