// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kL5pILS7VpiB4mDuhushSYLkVtgV6Ij+L4+ju7WPQeF6reFn4P0zdQpcdK8pOMO9NQBODwiDxW7h
JqS9o18CpuFufJGZ8IY3gcGc8IzKL+Ae8ah4YDTp0246AAWLKVEGS4dejqmzrRf/thXFQh+3whSh
P+NhMCLrO/I6JPU8X4xAktD8JcLpscmOo/1N/uOfriWBLQHfeLNlclz4bXx0fL4CBG426XcTZ+5m
1rHiWuUDUQOF1m5IBsZKjaqqsP+aJt0/tFQdmIFRvIfGBFrOJ/8G4A4myz7r2F2x2+nGFcT6J8OQ
aLiwW+j6gXRLEGNwbzrAEdHmn2LP3D76fQh6vg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
O3b43CJwwxNPFCI9NX21CIVhcOYoQpryiVdUZhijrM8L81HZgh/1bIExBQrsB9GqgvGAFrm/srAL
VLXbQhSqIcSyrS/mKMAzZV1HP23YZS1miA/pBgKiQmAt0qCkd8LaUD8Wk+cUHoeJat+gY1o62TUj
NTqSiHQtathg9X5f+QFB9550cBe5R/HUsILuGjClPLSPatQ0rf9HbjPSdGIzPeCYwEHQmGzrg9Dh
NXeCodq6c2SazZ2ReL8HLOeSf5VIHFZyTbJGs5lAdXH/WtVvVWfXCiiEMdM7YPy/O5JYtSSkUF7z
3RZxxT+5uiFPsktmTb8Eol6b0OejAHfOYADrgQ/bGeh50UC9WNLsdT+Mn2SP2go3Q5AhHCHnaSpe
pC18Wowj9djPzKkOFZcstziwyprkNLXbCgznAREZUhnisEEvGg7UvmyUBsR15LzX2YQY3n+6cbbC
PnLWay8t3PvuLWaVKCg84diBTeLdO04o/AXsN+NsTSmtl3PebPlmUqJ9nSdWeTFfDXat4hDR4WLG
WeanvSsmjJ1gijvWCAO1DnWtnnrq+XPMTgYsOPBNNza8bOsknlOR1r82xXfuVjF6Nlfi4Dl/CNnS
OBd4UV58s+WCODfD8BlLseuiKmBner3WsOmbI1CDxN3L3sfW3r+INdKaCy1W6pJf/oDX6qXSMfSM
1uQH+879LUGB8dWBO5MGM3yFY2RE0u0aJCHqj3I69j2UsRIdctFmYFDXZ3riBu+4Xu0Ii6xFJw/t
6/cM2AAJyKdpyao7fImmyuQ4PCRw9r/njCwP2R8Z5ef0by+7NXN/W/YQFgP81CX/TZNFUqlWypux
tfRalrfnmvYHkDOENeG/7/z9S09L52diytSt4VA/x9B6B4zsJaCC41Gihvy4Ip5pXYHsLEhrzhev
FRREodI6F/442Qk8OJWwcjZ+iXOtqw7ywN7vsGL+yD+oRekCW4I391RGfF2UBt69BMVU04a/Gfum
PXHEiDoKQvFJJJPDyBfQteDJLKFQ5CKRSKBo6e3piETxGlxuXo7B+AuSIwazXC5I5WLCe42cNmMa
DVRR/br1U6z67H3NPe5n1wouxB9d4MedryWypwlDEvLV99K8zYUfhZtcl3wq/JcYb3nzmNYwr7MA
WSHO7x29GUZ5OU+e6FConyBNUpLZgiqG20DDqoa0UrfAS7qFPgghB0fFAgA2NhBDhyUbqW9IZuR8
N8kNcCit8u9HhGQOxIE+dI3yHURq++kCpG7U0UCS7FyibHDfhZ3RQ2zV9qmKiNmR7v5WTlGhEGYK
rfA5ZxxaJef07W012MCtAz6s85dWlLPr2+5RVG06nJo3MZrQ7BLUdDEtbp+dZiQ3CgKjboGjw4QW
+FcwBpH0cIHhLq3ICaYZImfrXTzSJek+w4jq6n5BcD8aj+DZXCe6SkM6Y/tkJHmVefNayqT1HYM2
B1PEEQoSrqZgv51TgcloeLK32xpy63qmtdefnO5/nCJ0kjP2bCujK5Wxb6bTdaDv6OnIA1Ap8DtA
yRH5Jzh4brnOMJc5xDUw3sJZViVyCgenCAljQ7mpggTI9DUeLH8qziKTZI2ExJj3dDzuG4D4Nd7k
fDy7mwWdjxuIwkNtKh/U4tw5F+O3t98+0KMYlifw9F6wTfpBJeIMEeXJqX03HmL0CnrIkiMykCqh
IDqM/BLx3mJ28NWWotA/wP3q6062/5dV+ulzXncOqcRjA9AG1PyZdrsAVOYN3+sak8ZM7GN2NBYg
gRXhJ3Tei261guOr/zSxylcAfZxsYdiWSZnLIs+mdJojVM22PGasebQZwcKMs8CKAHNofgsrAtk6
+zl7cEq7rJvPaUhsVt6VWNgagaXkmSDMl3VxlbU5N/7kWhwXkgkFWJfTrGoB68rjw/eRyIZJHfMW
T/kQ/aamcqV8tiWET78/LkXz6wK2b9xNkMOxxaxYXY+qDb+aaKHC1zr1nd6sYDZj6hzoNmI2RCY1
sUbWYRSlD0r8+4RreiL/pVymapi7zob9RyEEEpM61f0Z/DakFhnnoYLqBH0NCGO4iyPOLz3b5I99
QjwrnVx+ategbe4yDCGYMF9FJ0KXy9YzvJ2sOXOlClKZyk7t19ltIVqtvX66MtHnsFQPiSQPyOgG
NPBMQMpNfZHsqFtksWLI1/1EpGgc7qQawYmTEp886I4PBVHLiGjkrd1qVQAfH75EdCqBKteWQnt9
b0BoKAfZsZ/0oBc+UI/Th8mIyVkKBr2aFt+yg6yq8RNkYvveSdUTeVR0ePKrxuNpECPXeWXcuCDF
t/fiGbL3Yc5gO1d/K9c3a4HeOO/j3LmqOJQS7ZN523cP+hQoTwLdtw3EMM2LmzNjQ5F1JZXcxTOp
GlBXRwrA4/DlCjNaOcEo/eXXZnhlGo6oQwK9iLmJir4hwzEqIpcl8ye+BlpVitSKJdkIYPAy99Wo
u/UcMuKev0pUUKg4Z55l+og437/aCAAocKlBwBTfr6NJ9+0/VI/o7PLcy7MS9Yy0j3vuFsm7GcH9
LHOG8F3d/cuY0TFTebslNIuOJABSp6cTdPw57BgxMcGP3cXpk7PAF8W4fRtaNUl6SHy2ku2zpP8P
RwZB6OEhu2Dz4RZLAvjneXHfJXkhjeyMZl5iEHng6rKIp12oR69dG1FQovGrAL9qGTMcMLhLvQ5U
vkOjfJBuNLZzaPE9UFa3ND/WzsB76kg7fH5XcIhn7MgIB8JAbK/hSRF3T2bgDsXzxddnr62DRila
SGm23zHD52r0qU/9cgSRuQZsfVF8BaryscivkGnwmlk8ulHUkAqPwkKQf/F2yDmGN9sqgyWbu7zZ
XpEtgo5gpJlZcFTOPbW8iin/xa47MPAPM/dAQWqlEDCle9aKKdGg+zWpQbhYSCksxwInjfe92syh
t0F1Gwr1SRowWaiPeRqnHjwS/bz373IkU/jXplh/5Bo0xaCxtVct+VEoLPLd7zcqN86wvtDr0AaG
9SPOMC55D+DpfhW8+Tn4ReHN3TrvPfsQl2IxQ42f1K7F+J2RMdSBP2iG7qveAOgHxHhMPnhxocj+
Iwj0VZlJUZp+Dzijy7o545/eW3QEgtK+YAxqDmWH5dLq0jbv9xe3XRpI5UQ94Cntd5qfuoEtJhg9
3nd/g7tzgxwRofw05t8wwZBZSImuniKkN5CJSZ3quPJdntdLR50GT/RsCux0ylA3clhLO0ElLJ6H
tVkxoyCyF4zxuoqimXKGF+K9s/Wzl4v1orjPcVs9GhsFk1G/0lJWMVZBLa4eL+GYgkmaWWuG+IUQ
upaeaoO1V0rzXVCB0V3L80G7Yu4hNEACNRS0u65EOJciktfh1/GdIpRxdKif5lQisYmstiDv1O/r
eAY3it++Do+p2sjqXHNBweD9DPnt4gt2ItaNQpCAHxJa3p+TGiqHNAHdsQ1R2rLY/glKVaDmP2jt
/KNkwYhoSFkQ2X4nuQOXsHoNwQeZMPjSIRt+ryyK+hnlCkb5Y1IQaUQfIynmkFrd7m2U25JZk8xg
bVBVhYsyEuAmShThu4FpDpo1eCZ/UkrBzYw5hA+HbnsQtPBUsc+teqEyUYUacaCFG50o3Wn3hvip
hIohikIFNpnLq7DbzFdyXStbk+amUXC/RyY7tg4r98kI2SjRBDd9hedvz1Qu6vDS3uGeEPR9wIrq
JKjiJZyI78QavyMqWlcsg0WIayD8RtvV5SEU6pU+UTNsHADtCAEAizt4pRlrzuG6iJ/AIBgUPFix
W2xeITiD5/RhEVmwGHPdygTYs2rfkgJI3zglDBCeGEoNcyPOKVHDBjla8E7rG38Ng9s1V7RayOvd
Tq2cov7w5o6zOEeZqulg5WJ1QDMi4tKD2JAMUFXt6NsQNac13e5uK3YRsOKPRXfB/ezZe5ycq8FE
xeWtBjXHr7j5CXiAfnwH3XuL4OyXM3ygHlkpNnbKfJ4U81/PjrBwUVck4jCyzgz39c9Bb8cucJ2T
ejvYKfeCXQxoHxAiI4A4+iBk6610khezOlUwAeog4uN+mMeutytGK7omjOC6Y7ZdqbOdlJCF+uW5
cSeKAUAnvSnnTSonGAhfFi+yN42iOZkU71leeF7/4RX4pjUTwoNVDuWdxLSjGPt6JQSihrlxxQca
Q3xC8Mr0RlV7bnD8LmSoimn2vWmlsXYu+/iYvynJ3r9DPBfD6XyBEfWfcdjpqQIFTdJ/gm7O8+Ko
geYnXjf1I7xiiIau1vvDiiYAEyI9HUcchED6ANyjpLU0d10B1O6BlgG9n/IdhLLEe6pcsuaRCOJ3
/PjLfeGtdVasSxtchb3ULH3rHOm9XYytHA/qd7DcXCrsjTv1D9S5XHj83/hcBsYbTpse1oGAriZd
9PjGHkMKaR2xVmOQLUIKmaG86Eea/LqHwVFwpoDAxqufb82+BOceeEvprXhFOcNvfnkkfNtx5s/9
xV32STbn8Ai1T7/zMfFxN6Uaw2RJljVTTKdHNRQIsmcsqus9+eGB1tLeQzZZv+pJiNtOppsUPNHT
hWL83MXunrJ6wPFQejROBk6IajtuqQtQwPv5FUDAEa2rnkAx5ZR67BV6O1GktOwGJveFzGagAz5D
FGssUDazGcESop5BxTKF19Hr2/q5DPSxyIVjjNb7oizmkfJ/KBvCR8n8qizZijQlDdfEDxPgSBVK
qdJPJQ/VK7/IvgiWiwqhmpO7mR7TPTNiEA+V5Ud3HQR8dcJHDwvz7bf6E7jNuo5wzzOoFcilbRSC
pqeQTv6ywM1T3CnugRkRL5/YTnZHAKjlrKs6gp780dRBHvqvTIDMJTRZMM8kGfB1pNnB+JJcffyj
7+x0tDFDL9WpB7xYkexsUzWVzJuSdwlAfixJNzslCJIrocgECohnQggCnzci6n+4Dpf1Mhv2n46j
dbIUQ6h8rKHjJpxZe3Dl89YYbTvBxrOOcTCcU+RDcIi48yOxl0pMSl/RJp4pmSk1+MuZ5yuQa9jO
04ttmT2X6oDN+1hfs1xsMK8o/i3lL/2opiFt7DxsI1IqM86OJ3bUv2TQiqua9ngovi8VQcDkN1FN
AILVLKAw9+UKBTFgTLrq4LQAE9Gw7Js1dxZPaz1IKN5XEvor//18+5TUSQ3ZsHUUSxADwA7lVJbg
XNCXEoZmiWZqhf/Lz6NH/TqZPauI0aaj7ewd/cZVRrOoS2WE2Z0HZ43xqvJFZbe0Bo64ZnF6xdpG
LFbi38kSjy5PEAvR7CgP/bJXGfvTn5xehOIPzgKOOMkvSqK6BOmFsP48NmsOqYGx2IB2HPW5KiNO
MisTRJFVtUsady3UUq0g734tYHRC6iFUFT//k+4WUu6mlrcS7owE+XNnuGT9qoQvQASgMA+Idthi
UplLudLMkpvLm3UY7BonXIvzK39YIsN8kUs0wE2gbuuwNbgiRq5oW/Pb+ntWVtAYe0b4u5hQ5RF/
IK0V25sX5cFFcOla3UFIq0Kz9DawWrEJtRk/pi4nlfgn8FqdvQjKqUWtnc81BVqfNRqkOF17TjCf
wgjrH+Nlf1p3zp6mvqldCAOTbbwo1pFD2MPmW0a0opBX33v0jI4hpUfel0ldEphWcQWEeZWS+Frm
Cck2k/ToU85/Fbm+VzB+Bn6qt+S/chfjetHYWhy583ws4bktG8dGrVY3Yc9CAHgzk85bpqO/WnPR
bgiRaU+MopA5OiAGa4xd6nxmERAcGKsF0PMNEfSjm6X9IDlqgUmDe89X4Zu0u6oLofuIKa31YmLN
IVAE5FRteXIlajBGpXr5U1jRuhLWSX2QpiCB5XoKeWP3yomii+K5vWMZVUCaBZ3mnb298zkMJXzl
9Db5S6zxKXY7inOY3wd7O/FmAPu0yh+xyEzxNkQxaaaHuNXRQkCIYkcUB15DhKplCNfrx/G1dyP6
hAQjY4z7y6wDJAzG/MgllzYv7eA6c9Wkddor/6e4wikzHK0hDIquxO95hVlxVVedlSYEbBhigSyr
Ktqm7NbBrrCQ+lFH9yQ4lGcxCdsff1RYxoekSHIhGDT6H0WfP3CtmzPVyBYIRvL1MG3Xq3HsfRhg
98sRCYo8W/13igVZedOiG3kPvwSiwn07z2U4Or+eyidYEaPwk/rpjLbCJp9Xo1m0pFrmQy+Fuf1v
HbG8kWxna+AzAxLvyQT3Uvcg2JABmN6oAicJ2+ougZPlNGoINYeVFBgWh+7g9NkjcQp/g+9X5AWA
jEI+sGgEANBhO5TSxdKuVwo6oGqe/8f1goAANe01LZR67vOE77cRjDum2EvafxlaFW+4JG91hQ8v
PvKCfon0wYqRUahfHkHhRHl/p/b4oS0JsG3n8y551WLN87UyBkPgNsJcO8z5mdCYz1mx273fIVIo
ACDWaRTgsyMJtGJPg401atu5a5h6V+H17hLFguUXPmtIVVQvRmG/8g0fDEWdWsCk2Y0ACNecX4m9
i9YNdmvjH92tfvWBvm8JAI+B+tj29/QCzSemBekdr0AboH0Zb7msHzbIuwPICG6L6WTA7haNFokz
Hgb3VGBIZJJz0/CUezFG0Ct8oei2jL7jXj6Oyqx45HhGSODXw4jMGmlSQpnnExfDCtQ1k1zfSOeT
yXpOKjug9lQIson9XTV/mF0UA1r3H0S5JyG+FTaBP3NOt534bui3u/7djQCOl+le17QeRG7oVTGD
K9d7CA78Y+I514NNzq4i+KN8fQkcXL8bzyRMknZNTwwTS90+tu7NiaPp0X1f6muVeJlv9CZRE1Fh
RdhsvpyXzdURS2ImuuaT/k6aQ+LvVy3uG5lLHLKhVWHka/OSHojtZOkVL0EqqWOEUZ4A4cknNRDF
cfTgOVHuHRVvyIGgatZKj9CqRUMYjklDWUhzurY8WjN4tIVVxH0ypmEMHjKR1BHzn+ErPGghVe9O
arbQn+gvhOKUYjbPq2NilCpUa5gktWQ/QtDxdiwS3w948/Ggw+iDQrShI/EXtnf1ZylLWKbI1xDG
s8c0Wdke5PcX/oN6ciIcmN0oXmAB/+GisCCkrWVbn7CGcalW0q3hiplUKudjfDwYsTDay9dcVpWp
BQXq5moExU666wveWEjrxMYJIqgSon6MDCcbGDDNAk5SUx5DdqJYbYpXSisX9r7X7iuA45FwFhVU
kni7p7kowQPFPvg8K9c8u3YiPXLRA9yOyay9Iz8sbz52E8oYUtv3HGxhIYNsqdxUOl4kGFQFqjVT
/VQdUFR4Xev1Giso/VbZIuAnoVweQ8A/ugun27JSmYkaFTfPxnYOUkMU0exKE5F0mJ3D9U+xuTJ9
3JKYXnIKLCR61ilmtnesYnuNoijhleJyeH7xkPWMUF36EIKkYPIEc8ikChMcDHFRA+ut24vKTYpc
tRI6RndCkDN/TKQQpD7QFX+cJX1wXvqN365GUWPBOsJ57LwBnvXxg8Hg1PWRyfjnuyUxSCuPQGsy
UCvm+4Zv52ZZXfo7YIXYVF69sVbLYTkmewoDUaJ64BOXKSykKAQk1vofq5b7OWeindASaVZEWWeW
CJdOF+YdFJ41siiBK1pVyEk1g0zg5fZ5TzpJRuQRGaS47ii9eVX4VRMCyrpT3OgueLoY9w9Hy3uG
HI5f6c+rVzvqf4es4hfyWNqVnf/htZzVl3ozB0kSxea3mJ3rpaUiIggS2Rd/zmMvTcXEqeVhYXo0
GWvjYP/U3WehbB6E9k56KXVyrj8pk9BtwdG/B74EWXY5S11nFwfPLkkoQYPTbvtyHXrjCsyM9S76
xcY6xTwlQbECAoA2cp/v0VMtLEr9N39kBthG74QCnE0VB3RPLmMnCiW6piXOC6IV1kVNNNb1ugy7
cX5k+eznTpUGXZvXBm00kpveoopHcCdPMZ8TZRRDAQi0dOSj5a+ylhNdbV7d3CXSnFubNt7OmKMZ
OFuVpAEdq2zp4xZVTRmJgu/J/nga75bFn8SOovoTx0bRqHiYWKRqzlBKNvjwM5DQDrOgdQMI5G2f
dx7Wrr9ciujV/CYdafDRfaw+ANk3OYs/rQyg8n1MmCQTCUxl6ChSLidDK7lKOuhivXXI3BRIcNNF
ZYWHzP0c3xdruw5dLBKdrXy62Pnd07CJuM9NsrHq307Osk0vJVuySfSlacbaI87cv+yZOBj2rvaf
hPC/g+1oTSwkd1Ak2aPA+Q6nI2gLNtbnHESG56E6YFoXpGmbXuqMD0Gv1Qn782maiz/vbCIBMW0/
cwbHQ+3xFq4m+PdNuyhYYieimsqPbUEUOENOpnnv3d2pEdRu1dL4KAZLYmcqW1g2uabIZ5sbCLvy
L75te5DVms7rWZJ2AClRbshwiQd6O7R4KvJedmvlUhE/1YTDbBVxFg7fG6uGETdN8EdCSvHF78wV
umd+6H+BmQRecZdISqi+MZCC9gDktY/DWNn8jMZVgDQJ/Gq99V6XuR08JkqIBUSO9Sz4FgnEMvK1
6BXQALuxRNX//lBKs+Gg6iOlNy1ggiODJcgGRew3QWUHdrcZp3pUkwR0FKYRg9rdK7gDgEjHzTT+
Zk/vfgi54uhnHnnmy2W8J+N5zdAqN/5FwzeQ4mmLja2she4rGEnGv1F2adOOl8dTy8C4ho+K9Fq1
pRcH+pYjgK0W2sjme2IDocm3gLtwGv9IR+hDyM3Ij9M87rriifDdjxD+iPJZRIpLh9yPylDLjrc2
moHz9uYJ7ZbAs5nJbmfq16DEVZWCPlqM/A+xzrqUDypoSPQaX5kdqZLwXF9pFgzQQDZEoQq9Bv54
t5f9oN2DvsW1sXiv1RQELrbav+t9nrWGW52Kv6IXvDImw4EbOceo9Pzj4FBwY1Bz9aTn1tILbiUz
+YiIEKb98FUgCos7Rju//c2SkUl+YcXSpd5juR/JZHLgKAJrKkyGEnbZabGlFjGH2Z6H9+vQkv7h
DiZFEWUYOZkcq892XhagF90DBWE6doPXYXFw8AxA58hMvXfcj9FgEWrWlxnFEE3EMO9Wl9mBe0an
D8GsJJZqXHm/wZkiUPcgD3ENxf1oZ4MMON3m8TrK4PckFMQstKxbG+tO86Sy6kxP1DLd9dVhM1Lg
IIqHe4+VqvmQlmm2jJ/X1FOnbTN/V2R2fYP66k+YgBe9rjUZ4iEwQoNBsYtCVKV34Vb6/OCjeRUj
a4PYkFfFSwPbhAi8X31+r8H+biAz85QvPXj4q7jO+H+XLwlk48xkICdi+HrAwWoF1pc43H8U3wPa
DVFwryQtq81GGnga3r8TquvifvEI3hsdI+DbKze9IQYB5RRjANCYHiOneC+kMZB7r5drk0GMZp/Y
5euQvLGW4MqNcep2lTN/BblKz/qALqmmUUPikH9TlVMmkIItL8zoEPcF4jFFrmI0fpnwN5jb1LKB
AyKbcu1XUP49s9AKsXO10rO1Efn3UwCaI5UgItC1oKmW41ZCnJwahnnCZ0eCSzCSHPuK9Fb0bZeL
HNpDeNUNyFN0oaP8HDhennU9BbLpDPKlqx5wJjBkJdjdf2+n2pvy/rlhVfw4XyvE7yAddJIsiB87
UWLM6b9asaXCt00NQrESpef5dXWOs81DEmQKR3wvw6+HfRD3UWxrhZcg57JY9mxlhl3wvIAzcDlQ
R4AEgknUeyvjPiLvm/YnnR8Z45v/xkE5rdT2sgXjf6BKEoawmwS+VAoUDaEvevPanbRFZYWzir90
F+s71gpRfMox/4Ncwznrfg6C/9eS+MyYh7Xgj+k3WpPK83w3YkdgDKvMcQu6jN6X7d3IABrsveYA
oOEpuQGnWnbc8Lk2x2zgT9IQxD1TLBage5lfwCAevjGDIiaPclmNrFjBLsv7gGguBbp9f/uBm7ZK
l2uVR7DHZuWMUUtWmNc3jnSX7qvcpw2Ktjo4xsBhtstHNHrLMkuIzCM0Y6Arv+6d5VFDvhsjyfCv
tecr3ecgXconcNv9fJEP75HWsI5PMCYlD/8krVQvXhe7u59ZYO9jR/oNcW3+oCeSI2X36XQsWfBA
C8GAjI2O6p7wQMU+kdT6qEpc6rlsclvpG2dzYHEhHSHt72AztCMCSiMU6/eTIFSVQB8d1r78KyTc
MHswV2VRWjhg5Q3zWUlx6nir79AXtpqKLEI9KgdCoDLJwnpNZ81/4gaR35hDEKRd5WXT2Mi5CR6J
2A2ZkrOQ4EZTVBOuZ92qcjtKMuKlSzwh6PRE/1kAWERXfSvZ49cOOQqwi5BtRxJqXM79WRKbmxVb
YLoRomiLlIzz4gOITf4f74EUsvBK+XrHCLyGPMBD42ydkLK0ozS+dz6+QorAZUIy3twIftQuyCQm
Iy49j0MhqC5p4Np65WXOTHBNgUmR+LCz0HoBy4eygVXeaZ+dtKWeF57oQSyv4B252urwUzmIAdUS
7uARuff/rGhYQR2Z2BIMbEpwnqb3r92QpPVlhZ26r2fna54eeYZjRy5O0ddnWahrEFbCSz3dNjji
5nBCVtSFAZcUrZloWSZdY75IO45gLGA3Sq9HiVZThPLyYCA9C4CV7FsLSzAbgc1VsYhvbajMVbRt
cVkBXXfx2pxGLkH7GQh0i+kp45399VhLbIsKJoWT0cT4LqQz5ZpDmq4rSJVA6FfNgvln+rkg9kdA
QNc8G5/Wffuah0odymCouALkAq7tiLWrn3sqYFYAH+aYOXG9xMlp65XEVuX56VnXzH0G53ZRrsqS
fvTZ8V5QtmduvKEQq1UWrlWo3UEnRDOy8tFGrEkCc8FryprHUi9ZiGmOT4xNoZi62ioRC8nK0pGe
KVohIU7px+iMHOW3qtaYbdsFNHWiiKIgCEc0rK+AzQ8K4QRoF81gsoOI4r+dxhJVU/l2452NUrOE
WwLwlpRdNBqCNzeCJiVb7b0GAoPuysYrhzdrmIAghlKcxZDZpV/xN2ozALvd2gWGMpuq/v4o6VgD
kiZrckPEMwfhGgVXMHkivNzMiTdt6oAxBdNxO/7OtoMF8wqC+Sfz1xCAsSVvYhkEOT9YHzCZ6ig6
yNjWjjuLqU4vqAEwBChmRDDn5Oouxixfd2b8Kygsl+wEd1VhDgatIvQ0/bXWZfZqLl4XixoC6dq2
D3NYnqZOcZmplwKQvY5nsxe5lUPsCSo96XDMUfOEMxvIdK1tCkKqYHADVyU76of2M/lXItMVlJ5J
4V1Aj7LqvBh/fB4naSlfzhcPtvak/HImqCemGlQXpyR0N8+yQdRdxPV5w5c99THrzu+q42LXOMqQ
PEh6h0VdEltqHufgo3uIF8DtOqWBU+jrY9GxKZb50RtcMEjVc8hl/7l3IchP3zKYzzxmvXkGQoeQ
EGaLoOqRrmaB8YMjyxnGgFZphOMSZ1/vKGU1eak+nFkmBPrdE7xdvBR501x9OAyHlHmFkJPyMbFP
HJP6C8vApUdddwlLP0SIEeYr2AJFq7tgPgL3jzRWCGjjk9EmTPzWL35hRXTJONlCo4744jxUgeKS
ZzJg8qySYR5RzPfAjBkuTGtGShriwR+yYxfUr0gkHHD/ptKpzXSB9dumxr4CAYQ2cSuyaETqbO6E
awBsLyCUYzIJthjtuabh1oy/VGQDe/CMG32CKUI7ooQBHyB1iN5sh/vH1SD/88B5Pbu7SOcHjtLG
RXdcj/Uyrzm6kqUV9l439Pifaeu3oFw/58T159TAGoxRgai5q8FuFQPwVh1UJ8oArlqT00q/gSFu
kv0pDZV27HnecsLfTP0YWfHgaO1HVpvdfsJknGCzkY2lfLjS49HobBAg+WxSyB257OB3dzZRBKjR
MWoRfUXcWk59r7VA1iwvpPpIF1A2fR2IOTOFL8ExO+XNjmH9ebFjLtOgEuxQ+zr2yaNob2lypeCt
lsEwihMw2BpDoLP45Ey3jA6a+SqPyEHgbQVunAuW59CYwcsGaSqNenc1Ps/eLCkwQ4/KOBVt53UV
darEdfhTrtTUEeNeO4MYBRreKTpxNKEP/WD2L/7AuVKMF1m81q2aSobxQ+D8ZKKbCXm1r+sg/LzH
Zjm4R0UXlwyKdo/b1jJOarWc8K4UqPWnhjU9Nno3iVSG6kcK0RreK+za4GOXELhlxPTX7SSPpl98
KyNqThKqJtnOtw++wZCI6isgAOavU0FAG3Lc0Vqx5m/Gia323PqwVuRPX+UECfD3UE46k1b4m7XM
FerJMdqJii5sy4Jiv9C1YagXsyzxz9OFGAFc2KkVD6KoFqdjLDERdef6mbVvJyERMKszYKSsjFHM
YZkocsDOeDC/IIy/XuEWaL0Chq5fQFC4gp1FeyIAmJ0KdIDLI2mbVAG/pu4BbNooprR2eoTr1Z6Y
AVvsJ4KnCNCavfiPixIwMfAmQBV4dG1JVhdugLbTrf+CXrDu2ONWVb3kYYGm+SJLaiCGR5a58+BK
uJ48OifG1+Ev6ZePi7bA/I3qr7K+w2Lj20vbOuCMDcmA7MV0MCHSK2v4uPVvhMlFqvpclQL7Dffx
HfB4Um6ORPFDkx5GK+lJ4sGbjC3Ld0BVzPVktWEcGot+bKFXl6GuA9caDcZ4qLSAaYJDk1f+d6sW
1B0een8vYvCUtDgFdhGa22gF0GBl0yj4/i9SmQa82bYCV8kq0Y5d1apRXs8iHxitKe9B8wtjtF3/
SWMqax2aStQm2VySqKUpeDSFZlzQ5aTHFbUp0OtLXARC6LreJuMvpBVa1Gfn7GNVuXDsGaaB7DKj
lo4JCG/K0Ifsuzz2t6kgMA9kBGgyDr6sv+mVjvjfvDUXHa2GKOmeKg7tysK9p0RgkVtuIXTViHU2
1AqdiPIJIHpVxf5W2ewjA49OkSj1zWA7pxxds4bnFSorf7Qqwb1+z/+JyOQyGxHBk/L9n3qKEQVO
i92uQ+bckPK8cj/XfZv7dRzsjnYcVh55PtR4yxo70dTJOeQhredgG/JFpxHABhhRyv2EwlL9dZAY
AxmtViXc7K7+eU4vXJFeg8NC+fcIKwpcgu8eN2TWeMIQWvUyBSeh1WepcAqkswDM420d12uVGR80
aRACM7eqRb5BA94PNVdIa+OGj9iqtwTGyEEHv449lXKEfpEEN4XrTgXJ0I69/YLf4KIyHmCGtqgO
umg5OmRjeJiOZekRz5LClWSxdT6WkRd3r0pH1eSsdxungvPeYqwQemwbUC7Vei2HGfKY/56VdTMO
HOXMiv8g6Tz4+R51hknYOVLrLJNPbMMxdD2BYmy1Dr8jFwJPyj24ElR6UwsE5N4yTXQ2MMrk2jB7
sUcqQVFIiqX+nNKQEA4npEZkrnnYP1Ha9vT0oaCBq7UIF9XbUZh18niu4WwkWYD4H0+8ECq5r7/F
YU/iek8vn9CqSa4YtQb+PhfoGtNmKrZx5CSCfeG6W3spi9vl+WNnp6fJVicSiuFhZ/eUsPt65NYQ
am5p05IGShaySr4zDJV+Qs6UuIgAjAnisP9kf2F7UwmIywO2ZwbSvS7c9kNCmYux1ahwnEH8hH6D
A2hnVFfbdoLzZqJir/3s84JZAIwkgQmeiZogp28HclfbmU6+sOOngx6A+U01OcVECfNRyrCZhYV0
v2qF1BPKUIg+vRVnPHQ6FEpz6W25IYVcvVzW7058A5QtSyMCCovylom+AfCQKrwRrZKv2lTZWrOu
w2FvSbS8d4cfP14HoZFfLCfZFoQ3MaynzdSwESmbyz/eM//oraPD5vLsPevFf+gr8vCgGI4u8HXR
L3tuWsE5IO9rZ32NgwEiiGXN8qPbDwe/krTXx5JDIT3QqUdMpsbsY/P95AkRZBvSiExhbfmKH0lM
YjI3DjPxnRJBz5iRZrvShwxNZPrhthZ7aJszX9wPXHym2DYj24kT+v7VU24HBGTQGVgqYXzvosLp
D/gECuJMiLda1vaJcANLT/tqzTJf66hFnzWseNpa8L7marrgBvBP7lfyFUxID7NUWmeQ5P0iQcIp
2ll8xvSNigMADzMu0Auify59MlC4up/LcpumWwfItIIfp9aRZiFj9vTnmsvydbQfFUA7cpdZlNrl
XwtsizBPHDy6ioMaWDffcr8MsXXou3FxRoRQRLnbx5fblxcM1ji9k0l+dkTrjxZpD9gcgtpkjgiA
k5nj+Y43SYN14pH5ZE8QbRpNqdtEaSE3VNRk0hwgGg4a4NRY4ZU65WVTV4KVuwVhkmE9UWyGEr7n
IabRGdMp6BXutA57o1IoDMjAyipXRWGNC70MY5pfObT6mv60Q4GZV4qNkVrbfgbv3YnRIYT1ebSW
/vgIcacQjJk5sIHTmTTgz47X3e6p1PwuNpxKpO1ufDwbMfiSGWbdO42hTBqX34+fQ1q6ySYL4una
XWllR1HoWs8aEpjr7Jm0MEwnQVUPKqfdNXys3IkQM9YAB+WuO9s1a4vKUXW7uKcnjRLlC2BZUzbG
dgls448JP8vdBmpSqxyrcZbucWQ6IXpvQg9WEroAVfDPkyOr5Ee138FTcF7lxsQFA7g2JS9mqgrN
m0dRsG9NghbKH++/ztU4EZi1SehWhWh0KBaAlYrhKxCHNkEPrbx4mQJeJ9dkBc1DDWvjBFVv9nCb
4c2/SHjAcs9/f0wTAjxk7IvifCftHABHwIPVD47bWiUZclXnROeYveYxfWOe0c/oueH+umLGV2HF
2ASnbg4ZcyB6Sy0zeEk2zRaS9jfYXecNhRxXZnVLu0dXeDPLV/kb61/HarkObpiP+XMiEA+b5NQz
qBMANwdQOViubYd3dj10gbXDcwTO5MEl9vp6GqnVyMbnboNmb1se5DKvxJLkzoIb0KhDy8v7pyRK
W2WF2EaupUU+gJ116LaSw44opJQ8ZJAMJtCocFqBKpdJrNZ4zd6W+Jf0GHnyzIbJ+nam6Hocpcw6
4iHCNiAXdqlL1/1tQFCtnS18z4rD1dn3M2TGiVko1soIdHJ4vnqEyOXmXRXrewxXhLrpwhASlFl7
5mZRkl/2Hi0ngeAeZDCclBbzTxu/aE4Hc4eNOHKtOMUEbZ+s81bC0rPgiwYt5Kw//FizyDXXeK+7
MxuTFfdyQdp2iCammycybJ2ri5p+0x/tFvEZgsgqY8VCA5KEPgPbWjE+ZsFKtw1oaiSrUQKEoomz
R2XoBz7krN8Lp7EkCNnYEBc4a2bQZX9hiE5SJHUMymxD/NGZ+v6CIBELbTdMMtzRuKBigK37tRkL
Iop0woYTIMiRAjJ5PAgq2vccHAGGmN2qW5wOLiwO4y6sa/0w5JtxaQp02Kte9Fpm58trRCH9lkzX
TvE2AKS9N/WFT00saEKUtBDOGNoWaOAXj9rjDxzuEmbHCqF/4ZwIQ/2ekALZNLC153quOam7T80/
ka71p764IHLQaAlfIWOfoYheUovsjXRhbouWqLXn3wXuzr9nX3V62NNFjSXNDoCv9osx2zjEetJx
3tzCaWGLBmiN5JWtpByu11ocZvF3QIII24GCPPRcFv9LVuoHbwNjeRTXxO8ac77p7D6KxRi2fGSH
Z39odSyJqB6E12RA1JpXUnXLBvYtPJKeEyCV8kByfsFGmt2bCbiyFo9K+TQ9jU+NV/Cn0FPyVwcY
NPOg3PYg78Ch6BXTVnqG0rw+4ELiMRwV/x9ip95871/OzSCRQCU0q1tFnvwL1YXBvaaglKwzXrtC
UbkNbAtezFSLmbrEnfxby+/c64w5V7SprlLQMzvmxAAar5po2bGrqdts2Dbz3ZkrALPuggfBHQKf
868mJFfHGFGuTEIR9eBDlN3bRIMvpYURfZVayKL8+ZWz6WnSLxgs39VPAk6LhN0lUZFQoQghDe89
ctK0jwRcTvb+XGgpoSdl4C4n7p6SNhFdZLMN+oZknwUVHsLLvw/o8oDIhRuCeg1rZ84319mTQrQX
r2c6oXeSkymbusrtRQlZxuTB78xaSu1Ea8SqqNK84/tnRXyv+mKHQDPaR+SJ5T4BpV4MCWsl9Rak
xK4T+4hmWAKmlbYSxEiPScc9w8wS+EFiVeYw4OSKUujbmEhF7Obsb1yuAefc8xNBeFspwBhYMOts
JwCh0ppskgvu1k1jsSj6UnbY44qwlP4Gu3S0f88QTiRsQ8FqHTFNL9hESExMcxUGlSKxqNDwBGtw
OWlWHHewnT9BN1HsXEYk78vTObQJNyOXwe79qDNfzQ0gAbTLbrXyzTagHQstrY2glbTfe0BSytzn
e9zbPeXvOAMMGCYb+C1DeMZj/6ahfDBXPYKl75iFO1Je+BsruU2yGDd2hc9dox81/7HShSuBQUOS
VT/T3dg/GisbrkuNPw12lnnIdlztRaBdIHSfyqescv96NO8u/b2+frhP3mNqLY222ArVxmNOw/JP
O3knpa0UvevgFSUkDp9ffiXrKwj19p9XRynLf9GQrWu8XKOhkJiFY9Q+XZTAvjDmiNLZ14Zyt81B
8E7aYW61GVyK32ZeZozV6VGMCfFDmQgZ0h2nZJi0ljOpsvQWWcAwSkYWnSkFIAJBG7JxgwAbLtki
dXj2ojE4+PC6I5uvHfQrA6yeuG0Tgh2262Lp8j9FHP6nYV+68exroFRcvwVqRyrnkk5zTvjHrO3X
PvDrd0em6RLlsGLNj/906fE+X3H43bz6R1+ZM9+++dV+oO+NJ1G79fE6WY4/0zA5cioxxhS2Cg3f
GtRpYeaVNtO3puJLx6dgg60EFM9njoj47n+uZmCkrqEsQd6xA6E/CqaJbUlilSSVjybKitpaF/Wh
W4SOII8t8EZURU3vqZeMEDvXk5ZT54v/0lRpMaBz+ef0PFdbU9JxkhhHrAjAYClDocfa8nkJ7MX5
twdnEJVRnchZz/JEf0qHXyszxqSqOzDugkPd1T5Wx4C64bxjJRzM4qAE50KAscPMG93d/Oln+xMr
3KsJsgiXISOD0S0Zwn+0ca6T5WUCycFbZCx/Ype2qrx+kNUeXf6vu1e9Ibseger6MUJ6kVMBKW1+
IInL4C3oDqbXI/iF7oBSLz52X9IoyiaqcV836a+Ii7CtAIoDy37VIADOEgKUt2P6z5jFbXLeaqm0
rWi4jskJ64Zbu1oPcsE1KxNBH3g8Qz4OAbn7OTha/8Fz7DYf+T1Ox0N6eN0cr5BNX/mPxWaXomOc
zoIBcNsN7arCb8LyTzPouBFdGoQDtWl9D94FvW1foFvYc+PasvPqaZ53FzjYVgxruFPjV0lYuL8l
MkPEUZUCbV9cLjFaPcMQHy8D9ev5JmVDvFmMW88MOmuh56zWsJor3pAxeVsgUMHQXHdIDg/s805W
0c372TU9uW/swYf7KcX+0kiJtQoyOnXh42C5eq76A2bGUn0z6uvQcekOUZPUs/aTFpqn2viKiGQ5
GnEOOW+IAaTyCa0GWN+QneqA01XLtqX9l8KWfbZaQ2D1Lt6VU8KeQXNnf553vv3ByyvxOLqewAvd
BZ6L1b7/iggaACu1aFHXn02aNgCYXKzTXo2zfMx+K4DhPdxUv3JI9ZfmJI1+/6omvzNo/bjZUpvb
DYM3oWvVgGkugr3gPAyC7YVKV1UHoaxf9FdywwkuR98ktOl8TqtHiRycYgo4kQd3uDNSR6SZ6oL8
83iMJUWa4bsY9G4+PmmwPBvMMKxQHsEvnRzrSymTYot7X4ztfroUeg9r1plKzuEGeZsfogrUZa0W
Hf9quBF/KjCfN2bWAGY8+Z0FeaOZddk/oxYZQu/eclWeAy9pg/xIw5ybf2+UV5Pk9GF1TuGHAvvg
X9pbGcs5czVsSMh6nSWKA/lGvTW1izscjtoLbM5e0GSxsKLB4HokD/zJdpba8jjVQQeelz4pRHaJ
+q7+LWC0jOye7bw2Op7n8DEKihY6C+2O/zW1bFpqpFtwfDuG3YRLocsOf7t6uc0aIyzpU4wxuxZG
eDQgqMMy0EO3yvqZpMHYmJ0KjxxW0yCo3ChqSO3iESb51EAtrhGGh79OQ2JJUAqAtH97lHQ/56Bn
6mHBDnM5TBRrGt+fhVhCdgL1Sr5+H+qh6zS6/WRkQ0JHsA+tW7QTAsPBz9SCvvn/ZEx8Jb9FtJof
1G+MH6LnFhxQ6AayP6j2yGqFUGAA76zScksi28X2irGbY70zhqulGu74jlk9IIOUFY5/oIQbEFPb
ZBg7rel/Pqy++6iaxYA/IpiCxufqov+RNK2jOsWEXlCk1LEnh5ohsZEcxJ1FduLJjdoO94hmr5UZ
A3KInP684/GH2cWy00PmKEoz1EJOz4c2awzglkCN1gMl1SOGN0xj0U45N71zisza4S0WtO7H4IyF
DH3MNAREc07iIXz1gk0hseJ2Yytt6iR5Q/35XY93y+pA35ARN9y0MeMmpTht9hGEmwW6ppMyqzH/
AOXAe7RV7m+HKrdrI++klXGu3UnaHzTYoCZj573vulJ/MVZqZGWl0nfUdZrbJJ28QwkzF4xG6yDt
iGbEmlIFBsHYaowOHDXeKNZS/HmL5J6DqUwTQf7j5sFEO3hGa3Fg0WfXdaYmNrQPIrAFJA3toOmg
liHI0tK1TSc3F3CjRisV+rhh8QPGeN52HLzhAxqMVja4CI0AeC7NERoX4ZNYzGl7RQgQdQi50oqm
cdonj0uFmMUgUyMFIJWV9gkGgvMtAiLoyl08nE/tb4aP7Aa3fMxqKPcxIwL9OKQ3mIpWomLmfRre
PWlXMowY49a16sEybPLkHE3q950SFGf9U+o0bzkMXNFItjxTZoh8FNanzIYSr4mcmqalVRBlYM+O
an30NG02j0KWCJiSO+bp0LS+Rb1vRX1+slLBduNMk/zRCAMfJ+kpyz+Ex4Jc5GvSEHqcLBjEliqK
8ZKEYQFY1ssFd+qUo+BCDriHZ7HcJl8QprH7k9I8JnFKDN5JQNxiUdWbFDaFeNs5OyJmPVrQtzRX
nLeHE7eZJhN1VwpD0CAoJ4Gcdn5TJg8D2/iAo3oZXEKuWQ61K/yOgZ7l89FXbABe+rL5SFR+10SZ
mcEhx5PHJn33qzFyRK1GOCEvdlIhr5fsK9krfHbzi234D8Z7tDCVHYrlzDYZlSEHPLMnBc6v55A/
x+svZa/o2fzkDv3ZdD3+LTJhjNvLg/LjXBFKUNvalCo3a/I7jlAuEa7Jg8pItvQfPwjCdsJZe4VH
fDz8G6v16pWeuxrsZzXmZ1Xu+1vYqDvxT3Qv8IzoQZmUf4IIRYKjsHK99GZXArtmO1DzCmX+OOBZ
TvE5idcANv+lIwuA0oAiqp9gSFTe/u0iMnBz2FpZGv9t9uNKs3i9PMbAPuF12VHbc5ZuiRA1ze87
MMd0jUmdddhuuc6L+TczMagdElVI3zstq5kRXfQXX8Z+mrvNmSNYkM25wtdhsR5TON+rO3re1toF
9e+eCnjeBPKf/JU8YypLEJNgl7/vbs+ZucB+TEfEYZCFm3FGYn3RkH3ZoqhhtC50CktAL9XNXCLo
dg0y8Yne57irV7qi7zVsb4a/kmMo1fbGbGCCt+gs27nptSqa30lcUlq6pULpssWsxBkd0OjWeBr6
8yZssWxEoKtJZnrdJ6r/LradwwwFp6gVlPlsaTT2Gcv/ahrliaM6xGHFKz4jL+nPSiN2VRJxZhgl
rM28JnLTVnYXFqRVW2F7eSKttmbGWYbi7xTkgUw1iMBXuQhFRL6PmWQcVFZCKZr+JKg0OUD/6NQD
hQvB/1EqnVjxVZixPAZ5QauytZU43ZO3xUcWFJ897ln9V1UGuOeeJ30kXOG+stzn9kD03wbLQicY
KLD4U+cHvqUhtae3oB7Sv18n+Go4cEybw7lHCNeuKSiW4vpvbSdoLZG+fpnwJElPyc8dWmua/KCS
IG7YAMq+bbX8uDoxB6fSFNhEgnGACMT/8pdJnyPEOBawm7l44glBqJ0SgELKKpVjO9dTuvdCQ8zZ
2EMcNwCQJX/iidIFiF6SxMkMMiVMamDHwjk/1XGDL4Pdl166QqWpVTM8RgdqBI13fJOa+u+bULGL
fkqg8WFruSPnrhj0yzCZqNoe33wydfYj6FdDIG9RWM8ujHcmNlvuryBaW1Pz2h2W4DwbiQZT7pRZ
YrPaQWogr7/xrVVAPRB5DComEtzOeCZKbBkaLzVjCGCY28afdqt0nIZfXPBt6l2zEnHkL5hQ6LwD
jFtlZijWP5BLsoZyVcTEU6Yp5PbabBz6T9h73TKGuW/SNk/FkrOP9NLnOjpNpclHKNx/XkN38pmw
uKjXi+QxZhVWuMp331uQM0PCjEbe60c63HqaXNFxGlkrt6Lf0rs0NSJAJL6JhPhqEfdPYRVhENxd
X10w/eAg1JYOk7EBlS9PQsbNQE9hwVxLZ0CqxrbXWVuPtTKMUN2/ILjCQHuneN36zNoSj4DbDzgS
gKtVC8ntwAQhYMY7Hy/XfXUWR8c5LteV2h7zS6geX9JmDwYqVt4rOnxOc0gfDXDq2SPNBbWPsebp
D5/YlxrCjIsnH50OWNrrgl2aRIZjm96WE+mG4Qfl5eLKN3GmKM2ykSRFyVEZ9GopYh5pbgr8iu6l
cyXt6Yz6ZvrokgBzUBuDhssdac07NYxw/EexP/qltkJ0G+0x9o8uEPk4g/Y77MK4WL7ZylX84RlK
hIp272zy7QLBbzHMr79uL9P9lKjhEfuim4q6RO8vzlYBqy21QN0qbQ7qerOMJYYR28ivjOFB47OU
nYEZ3o7tlKZp56HVI55gRy+7JffhnjEVhtp7383zZYa6H27crjcJyBz0lGJI3ijhVUU/R5HH0Pl0
GmcMibpBzWUyGRevLzqILFB43IuUNoswp50m9harjm6XnwrKb/aUQz3Zv1Uar3piQFOP1yf4ok+J
cRdwADgoOlyZ9s/rV5qpT3LLep9R8JC7hToN13yxWw+8lVJuuGVvCslWQt7zBzgAwkfH6GlmPXRk
FSbuES5HhHLOyQNykAlbZj56MH8n1hxIPb3zvmk12BwXxJGCLkEC1rWDmqnqremtQwTSvrp0lnCr
iiKXsROy6gTqSL3nIlSEoibjuvoBJiY5nNZLxpob1iDlAyl3526Alef0TNuWlSPCSBTGYzA6J5gO
FoC/2HcdO0yblt8E82wxBl8hSDGu8MFnRkWwoxdFnJZEpkTQyCrtgRf5vROzWIhjfVgEXt7u2uKc
yJAvLhX1HHJDdgI0Onkl4WATDImy3x0RdUc2Tbuvqhjt9d5qk6K2TwyfSM5Alrw2oIKGslmu10z6
JSV2xuZDipqCq5+5PE/clPRejALGk+5Xb1z6OnPEHiyj+ONMY4JlaiwypjzkPbLIp7J2umBmXYaY
RjsbLBcnGk4YBS1eDLM9KhihcFKPjRi0kjqcx2jF8UqHh3HbbqUnPLRx0OP13wx/CDQy5L5RcHIJ
SRpWNYOnUkS4XpceGvbQ6QWxv93kffEK41NWso7LdsJwm3Fw+W9pmU3edEX14WlKRrYQP1Ku9UTp
kB/ABhoZdfbFe2HO7Pp+XD0NeamqwczvmiKtF7MwofCXjHKBl+gdkPgfGLL0ZUyzwlLDvk3QBPaw
VPLgcDhtvPLd3gWpjuHkWuNmaruhGheUYO00mVpKo/uBWb/83dyIYepudJxgVRSS7MfsqVznRy/w
v3xSe0Pv1AGKGyM0r/nF71jlW32lwND8R+Ru+51z3WtwJ875JNqOnLQhr8jtoNpRtxAgK9PQqOmm
REI/OV5GAo4k+fXq96akb3H1ZW+sReF7NCzs4DklUuhJy+UQq8ul1QLNB2naTtkYj8q9ZHsATuKy
H4nG7KAKiSTkpTbHcm45V3jl3NVef/4Th8CUS6un0tTHsVDKG9BaUcsa8AG5o2kMA+bAfP5Rl6pB
yGBwNIUG450O/94Q0HQ8Il3Kuk6MkFO/3ILWFeatYqf39ZarDZ20a9PV4LdVY2ATzBrSq6vUy1yQ
KM63WsByBVkZhL9R/p30W3SeBIUcZDhodiNXDkmHlsLS7HCNP0ZGTMrsKt7YcM7GYNYhxhMyejah
+0DLrFf60GXn0uyZ0LcQ8MqoD/OFD8es1RAAAoV0QrJu2XO7Dc5iLmPSQDWFstTQXneNlu+9/l+b
E9zyWY9CdjGvLzA8FRR90TfVjpjMkLM7E9gjXDirlRswQIqIM6eIEk6+RpczX2qRLehYWLXBKDKb
lDHREQBM/G65hF8ZgrscYji07btapXN5358k+s6zq2EAR0V8a2lADFmecbC1rtKb/FaSZoofGDaX
CJ13qfU5phA/79lCG1DTzLrRipHTSaeybWLb+stGCz6tRB/6rwbfOJ4C28/U/DwOgrxBfFYs//JW
ThGSfzfw4fYbNL8dpvgxbpTiKGFke9UrkwnpsLbs14TnoaX+zJ4IuCAKGIwCXkHsh7wTk0B9eYkD
CF5J5PxL+Jmv5OOoRRfSNLOqv+KQ+XClKLRVBfr4wEPloKUSVTIFVRN7dM/AqoO4YxdoflTq3PPa
cZCr7Kzk7tyYrHc4ifppQTZFvi1JhBX4Q9VZM9ieijZ2P9eLQkZOXdgVopceE25dA5bQsufOnHAG
RRfi+uAFlnwNBSDbrAn5F3eQwFs6Nv8bTWPjLz3p++AAfDHw84Stj6RTbkQwsKO5wEkwB35Z2Yq7
lBsNJDpUHRSJEeIwCDSK4f3+Bvk8GUXtk9xKCB87tkN8TYrEIlvIYLZk0c01XNdr19ZSnuiC8G1X
qehOY6crlwZSdVJA/f/+ZXsjebr2+14ciuPv5Pz7tgMROrDcsr9n88Tkb935qDtvegkBOBvQJDNL
oK7hdGf6XA0j3hD0fxhNjDvxEceda6hrTuhQgtryP/xxZptoWTDawefTQbD5fVQogGLKc/vjAGxo
8QX07nkBNZn0XcAfqu90jco6V/Z09jhA0WkG4t4DTN7YCPU5NBa4DiT/CAPbuPl/e23sAQMb290J
ILIsMmEx3jkO5A/gKYdrC76oue7jqkp7DWXFGmptZmMdeulAywhRDt9YhIZgrn5f4j+9S0It5A1o
qqjlDPpTlbBK5HanCWxg8XYGOj64yxXC7LxvLHP8cJBzQu6gur5BaANeDXrjwPeIFK94P9DTgc5D
Eu4Jwtn1zc3hCFYVA5tPp1oEng0C2lemXfpEv/wOLTN4nrBkRyoQ3z/XU8PHkzqBTOrDZ2XcUb22
jayBLzIv1qn+zzWODImQOoXX9Rq+P7reeYKAfxPH7QlN70GhQQMJeBS5dJ9JqPOXSnU/Yl1fXuZ8
oTTONDuSbUWsmaHBug6ADNT17HO4fcLQU1czKacE5KWLgNe57EvDGgyACNV7z1Ua+xzjYZNfyIXo
XPdAegmKq2l63xJvLtElrVlW2YuOnq7rLvN6j93kYtp/g7gOrV7wesTSwFMdXGf+xTeo+XJDLPMT
NJIFOgr0hfiblSDgiMYwVe+5ysqiybxsUuFfkcxY6gYmAkMBaREoMn0yC9NAudKR9IfZAXEGGu0y
kHzGmJzfwwZZ1tZK2eXyi9/g2u8WcDUKLJyclL0g8UFCW6Nlt1ZABXjnY4FdDwpJIhvUL90cs8s2
i5wVkCsSOAUsjSWAJHpIqOQJst5KTOb6iYzbMTemH/hHX7G1zOBgmmEwuHwX8AApGdtV7BuKLm81
KQczgTV3lVuN4qmhvWXxGGIvRRXwVqld5LePr4PzmgfNtj5AoaEb4hJNOFSp+b9obstuR4dpYXqz
WLw5u+/1unhekRXNVlyopbHJtr2tKXopMXVMLSvV88GZ4lOdT74/YDf7uSgMzdQgFV4jn5j95ZLj
h63ZaL7QMcfNUUEMlMsgYDVjVMhRY9+5s6t7lNVGJ1++x50jIxxxeefTnbeQgtFQueA4PR6p8/v2
cONK+Q8CeJG7TANjKAiLg/UldKr84Ss3OAbPd5EY+IyLg4pxepbnMkd18ilf536Ivr97ijbBO5KC
nZIBtmyh9euJ32KzweMmD2vFdIiq6UsIgkDOY5zJ5RRmHoDzb2DV8O3W9/CwcfrKvK6oBYRE1UdP
9stjVV1DwixGWjeavnKnRPC958MqpauP9dAmeMLX1SUNQwc/EUJwF5wyGp8Xeks5PvZVk4qrb/ve
ztcKOeHc/a3WtDJiwr9R9MOvQk06GVUl2UPCyVagOiIaAYsQzLdb9aPeiykNFc2YE0zfQlqrOlUz
wMJMGG4OxyqV0Wt/N4KzxhNZC9sKPwuKQInE5qqLx0AJ1kkO98Ein0CHjZ/g0JgTIbBcIS0RR53g
87abdClBqy3bucr5cFbf5p03ExJig/38lzzTkv/auJrLQpP2hAlrhxnrM40RGtI+gDRs4VGFNRQ0
yFKXGZl9yMEIqsFRUcuKmNmZqsTAmy93V6Ye3Z0GGP3ZBGv+twbYkRRwZas0Fbl5zWd4yChU0o2/
I0+UV9iEvb8RhisV7VzbrTflpAQv2HNAc1sDEht2B9Nkv+Pjgm6fCpIBmsTOovgq8GDGMj04Ivey
QJOybQuQMR2taGaOylpbyIh9FStLF0G9BgsZHpLTS5heZ9f4ZUrSfMMDh9Q+Py+HiZ95YnyWx1Km
1lGiNBQKFFvXCcmbj0ivL2IG8UO37zgEBZ2D/BvRRUZR2+7MBQjT5+WXpMrzpIRX4+ouZdJstFpX
RoRjj2u4GBmEu0Vho47eanpBfNzeI5fBJUZqJdE2mP/7goiV0auKLKR0S46ONFpW2EBHbdmj6gCt
+1TM0+26U/EidN2nH3r8AHhbLjpYlvJJf+LjQUOoPA9NWireX013S8EeCR6UXxdMnE6FbKQXAz76
8eGFR4weeRWRbkjYvvxtb80sMZtwqxECaHKTtcFFsIvV1EK76WsJCrql427l3dNU2CrCAghgfyo8
Bbv4WFZY0LApzyVEMG+/cW+lH9NyquB/OvuW2meTZV4mDCmNzAnlLleN22EVi0GtMTUZdpU/G9lU
y84IesRv2+0X8qbtgK2spLbIQFee+SANAFpsh0xCgA3O/y+I9N4pzpFzTk245vYvK0EnZ41DKgjO
wSzpeyql2J8hd8qmn+FyssgshJD266rdLMRI3Ro447BfHfNAw8en+X/e7H+Pm79gYhCgJFKnQMpm
E8HK5H24y2NKJJ9lhkyKya+tFgdLFeDei3ZYJFumQRcbFw6vqpVfSmftQs38uExER646QQ4qOa+o
rKb+/AR012mKLlraJ6hrEortsys8PEJLeHA50evCKrFQENSgWHv4nhRneGC6uQa9bPrXjSRQxYZ9
0lL4gZfUw7YpR+QV+XU8VMg/tgWeqIeRXR2e/g+vAgj1F1V+Oul6jWEf894BzQdQJnmXkvulK5YM
DNKg0VBwDYWglCaR8EV+e/oEqDDqpz0taZu3xBzsua7l7CmgAUAZ/UJCMo26cIVdDlmWqcdnh+7X
6KELmkKBDq6VXNSpGBOO/xRzLUMcXpZvu0NuFCdxvngBEhICzlHivA9h1xTeEzRb+73z+7owo07V
7+ZiZurGOf+S1+Mm5qd19rExZNx3D0ApycuQMstkZ8UHM1aczBXoyDCaPRJoZQ+jUdeKu+Xw62zI
26FsK0SW2SNdXlmUf/9w+ny9O96mypPsXHHroePsZ3sngcAbcbi9HN0EbWMWj6To9L+ny2A6wiKO
+X8r+9XFpJ5t1zXEOM3/INA2Y1QG4LJ5e7JXex/gRhxn9Prg9NOGyBvXBox3RjiAuN0OFSb/Y1ci
Hc/bfp3YVQcjhqknVmFFqGUNOdg+vMgbBU/FgbzJHijVv+MFuTHs5BgoXGGTQ4c1Esa4kpxtDi/g
F+RAWUokInEZo7/tAcHUX1AsQMty21brMoZxJ1zF6pjJntDonGywjvUqxM4J5DIA6p9e563Jch2Q
aA+MyQ4k+QeX+iCuBFiXLFGa/4oZy7CdJNzqSQsp+8RV1ETuQ1kHhl3B/NdNXeRpVfHIUeXPhpk9
FHm6nkWyfmh6Y5Lq3cCI1tYcXiIO2lVlSW07fjs3q9ZZAMzTr0i2bhTRmSKS3M5/tzkzISd0bxZ2
ia38tXwsgng2/VInITeaumueTd5AFBdjkOMhy3b7w3dN5WvsrJ/F/0AoYEI/0BFjLPcEXI2Jegao
HSX+O3NS2/jpj9O6UrG0yfU0TbSZhRdLoWMgruOLgfRmSht3A+flHcyVnpg7A9DoOzLoWg4OFiaW
elzvY2gdvLZjb+K7O0k23YvhAWXOnYXjD0U4lz+zLIG1OhpMDl/R15UqgGPQtD7AaezuVJEwr6Eh
/IgRCDKwo/XBf0NXcvC7pPSaqHe4p8odeSMpoIscxuQ44CTA50cnRiAv+qbuguvFmBm1uElMzbBA
rKb/O46JzvT13rdcEYnNe6kjjA/3kfjjxqVH2zdPS1B9Vc211NWXyhmNsSnman2/KvtHrbTIl7NW
HxbZW7EXmT3BDfh07kOtdFU96CDB+Gf9zITsqB/iXUROqeo6/fK+zQQWjxpP/gVkmvdNOUPGPS6H
VL9wKr7c0n//E6ZJm7zyjtEaZfNue8jrc6zOpv7TEVUr85zBDMRezjSBvG4Rr5RY9jiDlEnAEvD0
ivoTbgjg67RoN9FLl4fRuVBCWO1xV6foojo8kx/eLnjIOCa4whjbMn4/x/xhN61qhLCTt5+aI8TD
cPBfnxO3adz3xJ5U2UnfNSvc3O6pgTwapMjaQUZBOou0uEbqP6VfEnT3QaZknD0rjvGcRBwKbX91
nhNAzgd+azzI4YL56nGUO5UJTlQyIXxX1cJRX2OBoigqexqGOFttrpUHs+60srR6RYQEdR8eQPQb
Ho/xpPDFaFkj2/6y2BnwdN4M5KDJRmivLorRMlBzmQtNNVWGfSxYognW0W1FAuhiXqyivrNvY/sl
7rMQVf74WcriXe0ZVyF1uQFHo/MOuzl8Y7bQdDzLpEH46Ocz5G2s6ngromu/2I21hJ9w1rnHIaP+
nmUcYdwO68T7VirdtMCo8fceTDYnuMoN6pmk6edJc8xQiiUlDtQPbse2wDrJLvnjt50ic64rAI7O
4PDU3vC6v5+7zSi+Z7FfqxbqLxp6ihBqkMBXGuCehGlhZNnLIC889Kd7WK+9lEPRxCXRqNAvpze6
e5SlkCNx7Y3cb4WL47RZUEk73pFjftWmLiHlFhiyLjZ4V77FqvSqgYjncDCxmGXKqeLN6ymbMHxE
Ejvf0Vb4R8jCL+73DFqf1PByRodS2xLz6rpE39T+FQ57QIJui+KDP6l+btR7dSgXPXKwXrT+a18y
w9mEm/S9ADafEgMzwMoM89dTvd8Qr0kLBz6ehkQmBiRCifOJbFvXL1XnVaziGDE35laBbV0AX/Si
HunJ6goooStJ5nZgvduYtmPvKpAZBhRVvJZl9koWrK2Gmu9L0Nd16DcuVH1BIIPUGdhYVoBPeJ9o
dbaYEtXBV2OcuY7j2kjeT9r2z7ZHFzjMRd1PvfAuKOdhZb8z3pJrDCSQSfiso/3BZIyXepd/ljTU
fMFXAG19AFDD2PbOGnG/YRg09ubKjo0FBxNiYbDo5PlIWEbW7+d5bTuSgPCX5rCe9GigZ56NrJ2a
7pS2RzWd8hlDEpO91icCbcloxDtq/K2r59QEPt6d5abSefrzJkIdp589fEG25S8t4TduCzLVNkaC
LNaSNtenBZo4GBdFimjQIMAlmwbJ7NWl/bq3DH6G7S1elPUVKDwCCdM4ghxyfeYlU3LI75lrKuuS
qiTsgcAvZ5ZZY0VOa0vEjWUgzjUJpCYufqXrTwkJqgG5B3R7PIiFNAQQA7UiqujIFYwG0Qv13B5u
PQbINWuwaEFewTLYeHr1vS7dJPqJU6JI3OAi0K6/zxq0zyPhfU0z0TRPF73wYmp++bsqXKOVm9q1
/xFToZxQHa4G7dhIuBi+u/xugRCpnxsfsU8CA5S8uRtlhaGMNuq2Z+gZqf2NAmjAOlK8nbUEZAms
gfTXsODS6gBVCWmrXWDrd2WehEeBrG/fxk2TEYc5B2MVcQSRj5UB9Q0HlBh8PAs1DWnDfsKMKZaK
2woSMdEQlZ64Xc2ilVC+15yn1wHuvewtZgacHW4wsfhhv6i0OTG8eyXVuvggT/tMwX5QrzDXr/j+
pD37Wqzrqd7ttIIepSE6RnGytir9ig3hUa7F7VEzy+SaKwKqEvYFSo5ick42J4fqbaajLQUNtTeg
CtwNwyu8KPhadChporIBRQkVdaFri9CsVifNXU9LE2VWEae57vNyNykYUCnD5X8aBmT64t7Tj+Bq
p1oWGw3yvam2lUCZ1WRzRxaSw8IipW+cKhaetwyPaI90m5ovRLHBI3h5n37PDdyzsg/cnoDlP9NF
SNePKXIzCPlRr1yvxVQpFwyYgFVuJJOyIWef1PGk84cDTwt4CN620T3Jk743qDLZDYTTW04nG8yE
YDb12QwsIfjQWiJkmy9bYEATF+flVE+lMwzQxAZOZAs3jPC4t9xXuc82MnOD/f/NKffLjaFfWhZh
YfNY7VVXU4JA6MF9RpyAI4026YGVQH6o/odffLh+ew9V6yGXPGw3YkeclEmfcG9fkLAPR3ADNeeg
iebgjK2t6mUo00HS0n6EmYtNUtObgIhYECc6MWJUq2C64QZdV2Qx2n5EE1R74+9Krw0q5BjYBpei
EdXYv0M/C5+RSLb4uHSVx+XvZ/57zXjoqtn+asHosxwNoaleZvwcfgGIvtL5ecdXzUvjmL97/v9H
k/6GL/iWY5K90M51EA7Y2PTaDYVB3Qbj+UNlNDIqHf4MN9ZnUUYvxe9B/MrrN3IGHs+YBk3E5Wpp
Gu885D9rXYA9pz0J7Z8V/9kizufmprwTljUUOFGVfaTPaRWDYCwsj242xOXGeIzQceitJru0FTpK
OmSjIQ5qOij0Ra9Wk27RGkAz9dJeE50qhano4DZAix7en1jalnvz+Qqq7774aP6tuEMG33l4P6rK
3HX2GYj9N0EeAa1KE6CQrBLgvtm0SeFtqx/mVHHVY9HTLat3GkY1UHLbFPUnjqmxReMsE8DlIf+0
8Ujhs8ZxLK5vjcInjcsSoSxeqxG4VzYamBhVhpSO2cCerC1ONZ/QrBCYD2CgKF/PHJzHxE7UzHQW
xUWJZpgE1k00g84YPNs4tFW7m1PsovIYFcM6SbBsQlvSzxXHunP1EWF7t4bKWUabYWknnwBnd9+i
T6WDhkqR9a4qdJ/h+PjxwhDY+aK9WjovMOdWadOFidSJfsXZv2Zr7O+AGHmUx5pX884OLv1QK3qT
10rEFw/4szkjxsDnJt0FvpFI0GOf26VRy0b1tsMjFON08fsx/HuwX/51gpsfKEnv49seCzgCb0ym
getL7YsHVGYjRZJtJsT3pdNzOwuLVV+Krbfl2pMO9myi952ePD6+SR2yAnnCaBR8gukSASRO1+Jo
jOxfrt00QQy0RiYYwjUMpwpJCNdEj3Sz804AYxT7gjgCUsiGqQK5lE9rqTg6nbqgCMgFhr3TLGvW
uqNN0S8rPssEXN4xDQ4mIzbvdT7vrQPgvn02nt9ak+DRI+HIc+05BorybEKEUuvBM/3Tne1hXVjM
Lu85xGjllAI34SubIXsFvx9wJcAJZ9XltCNdAq2lFzqQGoO5Z9DZ+sHiDNvh3OAQtF4l79i9uJZZ
yahRVGUD+XxUCdtk6bBN7tdzV2yLMtXVPA1+gOooqxQAsdr+DY9BqzbuugTfxOIC6ujIyy3K9Jea
h1/KPd/YWx03Ix9Or74IwyElsgYMpMzhTfvKQI6G0n5oPMYqaAyYoL2gzgRRO3yiRtP9a0iXKecU
E4L57O75IbHZxFi5kbKkt0QgP06EHDGhe09X+QfAPU5zer9GtFD3yooYmIGIkLZc7VQgwwx2TXZ/
IBOpIZu4gxqeI/ChwYMXbL4ueUdu8X9NBygZ7pgD/Ec3UAh1ZyHB2a3Zlos/wByhMd8a9lmjOCx+
ORvDj+imUYLnrTRLtT/10kESnKDKwlnGscd06NxkzOBtw96LUDsHnQ15JJh0zROGjDGaFOvWyq9p
ijM7I422aEMxQXfFZIHguVkmjV1JU07+vXzhPyAQIqOH47yEVG+AyrYiUZeIyyE7ZVI76V5Bh7mH
6/mlIfTb2LZjo8XmjO1CPyJZ+kkxHNL3bZ16lk+EcYOfDigvjIl+vgo2FwTQBLv+HkPDngGr0dvD
VYNUKCwM/Qm6BdUKtQ432pEqw6SzttgSkFgY8NPsjR01qHk531m86n1YxWmiDOJNTXEf7R2EFsPZ
zB1kYPVj+z5HdZLjxZLqaoDdGug4CwL2bfnPqbtypqBek66wyVrvemeYEVrltS1H/Byl0Vm4t8KT
+zoEtMUdGpbgObikCGZZn/LgU8C/O9ECJ/0qDjh1p3onZwfuZIDY8NoCDMPRwHoTITN+0euuPKJZ
VQoaC5Kxl9vEBOztd0AvWUD4yWVIYz4CeqXAuKDPXffrreyHbKPy8siZAd26kLQlxMBb8lHMqodU
Hg6qCcWESlLzt7TNE+3RaAwntp+lQFfDPvQWmRrHfHGvnluab4/HzjCPaqd6VdjP6eNGcNJf92PW
QIx3+d9p73tY6KTWmJxfPP96hdcJf2KC1V/gy9wG/jl/65WOu6Ip9IBBZ9OJOZQ1PVMCsAYCTPFj
WCrsyPbEATmcRK9PF8ClJ9devyOTvgokq5tSqb6w1rmnqggK8dBs3Ttj/1Udz0cwZ7ZV1/vN7G83
Ez2DJGmbYt+eZGt+/M+RvU0B5pWCiqwMlIO/GJSLzglTIudeDvaFFfnODqprZ0JCXAwPdWmEa9KU
vkIc/0tgYvf0L/+zE1pA0SJthm1TC5T2YphMiRkRL0KFLgtBwR+ZV0AABk7FVX0koX4o3N04uaWx
bvr9huF9Gui8AtaHWh2vRNPHdfXJNscsSnLKNohzoyfAVU8eAJul9/QsHuMcZRQP4ZSOa6d5Kdzp
3U1hqA9PI/GGFYfLlTU+s9sXqQJ1JtUbvlogfiorBSW3oaqvZSZ45rxJEhXCZzd1N6aTwGBg9+n/
YU/87yHIXU2qSPPvMUYbf37qPX4B9olVVvOUVM5U4GPoi+XJrOQTe0F7+/vIyziZ9xiJ2kvJJgH9
t/R+gA7NpOKoM2PoIq516BdigwLt5yJVWfGave3yTucPzToBdojo1MsHANYEfhB5z21bkHqXxCx6
bkuw+Fqwn7VaFbubzxSWwifKX21yo+Ow6J2KUPp4zNP/CwAw2pUthy+gL2rz1W36rVQ9HGp3wYLO
e3KkiqGk7uWJ3Darl7pM5QgQWfkSqR2uxc5dMQLpyCUy8LaUgpEpBlMo2uvIgN/o/1TFvCrr70Nb
QPTS9SifJrbLerpxMw/PkFlxD1As8cYCqEysPQFlqqP2dKhnPvpBrqQY/xRNrc01PdW81rYBNBKx
0pmzlHmGTU+8jTND5OtRIG/vB54SyMCr9ZFO7mlAMf49FlfRT5DWlm3ct4V6xjMe0fGM1G7GbBEh
kabZTh9qWwr46ScE3v9jo3LDQB/9TZJw1IbWlltWHfhf1M42BhAJAa7erUP8ZA1NTD3XQUskCnCT
u01uFE6aUd6a+NvXjVJQmijwmbyqFh0JOZISS5Nzrv2LKuo3ye5GGESzF/OYRT2w1IX2PZNS89/G
hqazCwPxk9vSKSNkzgPvk9tY7Wjsz6zEe9oCQd6BPJOdDAYMmDyjIZyNABzlyV8tRzvEAZ5tvLY+
T8YUNsrTXTc4XK8iS5ERNyqdyYHE2/7aBda0bMjrMgmVlFi1NTVVG4pFLp29Ri7aggUGoCBpbFD3
EJE2HaUWaesHfI8eGLObepyvE8nrHQAb81PeFrS7+tyEk+XlWfSIXcSdyy/tiby79DLoZWg0YDtv
FVXOQuI8AEPNEuI14TAGbCikFFgl9R3xOLP3+QdiHfD30n7kZ1eCds476MhsVUxx+VSqRKm1jGc+
XzZoVosjRbkdlSA0mSYfOGMGsQekFpBmHnRWm16u497jlpMSnG2BnbexehfK8PkBsOVuhOaHGjdX
rePNavU1bATFbbUr+JwKrP/rW3IFR2xIQumTJDKQZwMKn4OrBrEpjiV20HvQicg9mvQqVRFz+79W
s/W1HfpVml4ab3iW+vyeAMy50CYsdz1pgXau6D8+4efCSNqzZBOVk7eTjP6bZkcC3c+XTfAiOPFe
NjSglbCmsauLIp7ZBVgohPBFclJ3YECgkXXhdFCyOOL3UMKnenvRErsXL4lFoPyruMSIjykFpQno
5OETCjwmolfXdpBKJW9ppjzxuAu6Rfzs1YOUyPJtpBW5pJRdKRVYGCmZ4jZo9WaB5U6nDdxq9jsw
79FjG41Z+USFW7TSnwpmd4iRQa0WbHwF4MmcUjKFnFW71JtCc406oOQVHZigXQwnvG9dtKaF4rHf
pBXRMRyjTdWL80WNM7lzkY/Eqv3R85MBpbjk9IBuK8/jCTFwpcNK3Bojp45AWd52TJr2/xgtIxCL
8zv+bpyaKHv5CY+XgSYDPYH+aY8Wiikhq9SPTPsw+Rzlsi4cligdBKHxGUPH4j2lOuAdRhaGTJoF
VEFAsZXiKxt6AE9KBqtc6xC8JDiEaxY7hq9kLsnyEkllWtKdL03tIQwOoo5p03FNw607VnQVVRaT
sMWcOD0oqQr0kX4dQSwW9Bm5QbafIj8e8Mc7V1HOik+suuTqjwVPgVWEtIK+Q3w8UuGwp0FJPVbR
xjnMUM5y1fI0fGFRhRtzhbQDfMz/LL3ZMGgJFrQy+BVpS9pVNwyU5npueIW9W4jZ41kiGgtl4f7r
KL60pNGru5CYBFgHGqHNmS6Pzn250zx986IwURFz2hgPsFW/Auy9dlYYJS3vgxWV2IuCUOX1+O6z
EvMFjgp/7SgvYmWbFZLDjl/Dtz7+qRXnaeopqtKWxnCks6tX8fzwUkxgFKAhyg4AzwxwjQJ63fCM
POxlWSTIiAkDwMdTGPl7LyOxr/fTfihmvpZua3Y8Dh5Uzyb0Gc0XL8qzHnrgVVb+oUs+eWsSh+Wt
gXVHezzDStGPjYOAK2500bGhu0E4qMKaSNdA31Z10TRoTf5W
`pragma protect end_protected
