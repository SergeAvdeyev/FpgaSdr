// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zv0c0zSsn34rer/QMLW6N4gfCtoGKxzquXDGACgK77YeUWKAtbHzO84i2JYxL17k
rZJHcD6hAi/yQkXeMyGoXq0USvlVPD/vZn10DZW/ALAqqPlIiSQR6PszwuP8Uve7
NcXkUCVgskYQwnzXQ6GuEjk0xsz6tFABjFKP3s7ji3o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
6UUicqQODZZ11f0mn/fLTWpv4j+LSWU86SqSQO2I+H/Vi3zhbqolV5nYpnV4szho
Ief3wRESYMy7doUfLJg9Hu43MWuH2eSCW/rnUc2Jlxia7cxTe/vNmC82INMAg0tn
8RMR7ZQJvN0Yw5qB6UEnKsICc5XAmzbMhx0DjnfxAsOmkM53leYH5MeY/gPKhdqj
6xmdfzlPKVbt1tjp6MjdXLSUkGhjg6n7E5DPszz1c84kFNVXUH712p/fW09nwS/i
tGubDOnzW9SCZ1sb2gtfqAHxo2KV0Xo1Tafqny7kWIrEaArusURn5uJX7mbFbEIC
qeT3ZUYcg0Zo57lgHWcqyBaPedpMj53aa92tIQCS7V5sEqu2WSkVka9EcjVtfO6n
RXNe1X9KZrgkoeodfEypXrU87LUay6WlKCYu4AfWu1VxOcZaCw5ZISGAgf5qHyj3
cFlCooCEHfPEwAGYa1hehO48kX8TglJBwiuw87Rtecbdv9LGRoTNNsrmgKp73wIX
HoGwY9KL5deQ7hhrFAPxAwW0yX3TZPTaKZp4y4UOvZeVCEY29oMQoU0dD7i53roS
6viOSSSZyZIqKVi/5NZEmCyMaU5uGC+BIkiYZs/FjjlOWEVZTDtz3SLbQxgXO52V
VHLY1ZrqiScOEASN5Y9PyR3Tol33l8CQXfv6hd7nln527IbzE5a3UvdMgvVViFeI
Zg/+xF4KPplCoK368G4M2DzvYb99Wf7YXmE86R4oRvGS5NDGD0Of+yOvuXknkixz
bbL14t7LsZHIKfMWi/nUe+Xp1IMoIoyfFuLDDrAls28VVVriQbb4Pe9MAVzsOIHn
xmE4x47rttavtpBzSkcvBoExvUOPkAx6BMa6bvSRE/FqyVDSR7CIC0VawZxm8sA/
a8j6ErNN0SwyqrgEseAD2Pxa4nh0YsloRMQmTRSjaKqvysiY6xTHeKhXn9tIG3gd
nAE2atfbjAbXXd+Ew6R458NOJXhoGqv0VS7Z8z/rOFqzM5WBW4ELZSaIOzcNMguG
iPGLapQojib956XWD6FNHagfBNJPwgGoSG/5oiciKb79Kaca/TLEddakam6V+jcL
Uz40rlIXryCLQq3m5DZDkzgnN5q1dmuJi16SfFeQtT2jcJSXAIM6jZkGud2tJrLP
FRuOnoc5DZHWiVNQuSsNpX/U/N6AKJftagenE52HVHl7KSsqI6tV5U3afev7M48j
aymBfCK1NH5zf+ZNQ5yEOzgeOtHZneH9UhnaQvj2PAU6Wtt4pYyqY7Souxy2K1VL
DiJMsdgUKV734vN/c7vJ7vjb+67w7VaZAMczlINMvCGUpM05rCFCQrN4h6ltVCzG
tD4kUh5DU8rdsDm/C5k6mu8ThKtSwsN0PtRZUFnz/Z+ZJM3TFQg1V14ZC3iQOKLW
qsrrfDEORloN7ReEY+d/Kh1pUmV2NnRweB59C912EqoN8hTcZZ9secP5/JI5GC+0
VkZak9GaRHX6Bolkm0bqI2VSJMI9oCzOcZ8+aA5mmqTIsk1R3YxlzV/oqpErz6wb
Ni36BwxE9PlnQGWZRNvXHSAiyhopzsgqw6fQ8eXfwH9fJ4fFwJsJ8mKil5pjGwSM
3V5LgP7xd9AAmQOoSpa1FJoLHgRLMTBVT3t6PsGw09xsKkKJii4/E5ls1p4isFDc
rN+Ztrj+WhYkSAePWWbgwloi9A3qoG1z6zsX7m07b2Drvd/+k7NboT9XsG6UGwKF
pbrOd/Zhd7vKoB74GmsXv0eBkAZKdtaRAN+gSv76AAIFDsDl3luV9m1YOffzgPIm
vnd2c+D4YiSaMS6550qBOmI2mGMTS/s808uK1RaWWYrxPVF2fTjR+gMQAQyNW284
HswcuLP5pQE0gkHnqABI1LBWr1HZasGhA4YOphMqmzj5uQsSSd71Aeo69epFG9HQ
YihGFNgmWIuQXjl+sfgKOKjDhQLf7dqqV8jOksjFwUea47HJN2186hX0F7Tbhu2A
hdwLtqS0P7Tzro8yli8xucQ6cXgVZ+nwK7Xp7rxtXdmBXSMI/rz9D4aWWCCFZ+uP
EaccRW5+0fof3Y8PqcOaeDI79n4H27hiX1jBsB5Bl3lUeaweNu2GkXLQJjQkRTFX
2lCD28hlmlT8ST6PJ3wZqKfD5PKk7NW6C2X5RF1B8HDjrX2bkymm+zep6vfQ0wo0
cpeM8I6R7Echukk6XCYCkbBjy+vrmIAlHNB6dQzQPS38FDu9QD+854m8aYi6TNm3
o7tyi6Ixxxt8XxUCLrp0+bZZPzNxrbfGPGlUUO+7ajGNRz8U2E+qRNjsSSF7Caux
MOkJV9DawxfnKfsoRtnYazY+UKuPOt5ouJHI1p0cGLix73IKKc5/Z+AIx0ChEF20
6iJPoHA3UA2DyCD1ZO4HIhEzBEtUzg/SsT3uD1G+eppjZnru9qaIIWdVyqiqqZ2s
CRVgJfljntzPtbjz9WJU1OLaOZYkBwk0gOE8+KAZNFv2RdN2vk1v6pSR72DpBSm1
5BsxjwAu5konrQ7P0kCmmRWrJdxG7k4WzLQYwFTlgelt4bx0v6tu6TYeitp7aCBR
pFzkqC9cdU1DH8OTO66OMjjs0UJT3wIrE+ljyBjBnAcfdVO9AwtAADBoGl5OWyQS
CHLLqiKahod+TdrGFG6WQZi26BkNK4bjJn4PfwRl+9/ahaSQ+L50ZN2SWXDpBOIi
dyrxktsKhj3xIWrA0q/D5sF37nBKtLm1cS+EtR0GjXcJ88ol7ABHUkXD3XDpwUpO
T/M3iwHkgDG9oXLLRb8ZNB3njz4WRP6AqyleMduXRA9kJJaHfZm7wCyRFxG/CDsV
KItjNS1Oxl7fGN2UastDdUlphvPEV7D1MD9Z4GCSCKwXGAWBDT0JxFf8w5K5RHzT
oWh3FCk+NtwS1BsFw7D2LZZEdzRCCfUFmeN67EefQYfhFcLD1i+oLHeSwwpXGFst
b/zRlTQLvm/JlmcKMTyNKdiGpaRTH4UDijIsIc0T2zFeEc20sILlvAK2bpWhkNfn
lAnFltqFviRDR8Ve7B69E8SosfH2bAfS6Wo5LkzC1Pi2F86Q0HQsa+J4Spz/ZDko
fI3y92ROjRZGkT8BgGGyu95DdAO1dVAmRiTqP1kdGx7pnAWw13rg7ZhzR2QDYF+t
SkEPbesszAFrVEZjTZwnyRjRtG4bwfF7oAl3z4be8g3fIaXeN2+o2ataGfy/De6y
zKukPp3mTkDpYspOH8TIl18IoIkMA0MALN6P/9FMhZftjVCtiMOAW93+U6fkMhWj
+JmwxWfVsNGWKzU4GQo0wVi8cVyxi5fGS43dxmXwa0yCnH2tic54e8KJXV7yTSak
fhLC+miF5E7CSnUlmfCzuZpxZZm2m96ACtxO+lUo0J/S3pGYfnHVYCwjuMcqwViz
eg7TspIiKB6LFi0uz/KmVayyGfP02LtsYeSkdLrui/oQ78+4eBHTwWYiH8XW5qp8
pDyPz9KnFzLmOf3B1hi5Es19mARxdWN+LJUBSH6KsOb+QTibwMz5ZbsP5BsLyn+P
/Cmh9EpS840v/yJKNZ265615LNa6SbflbE3lrRZnknbsWQtlYaGG4DNt9x5hFGj/
orXQaPgbtlmmh4G9OxOf+LOsQN9ViBCPIiZqcm4uPhO+jZwm923DsqTVBR1EeUI3
D717jIy/j66nSHefHlrC5ww0CvVCiB7PKw7vyH1pfNhyoMFo1o/xdpwmJIRwkD6p
fkRZkOGBkZiLd30ZQnrGFzGoL4Ou7bWJFdUYbfkuVfcN2q1NdDM934E0MJSsRvi8
TvH/iYLz6tcH7xPAFfVeOcmi44xD49SPF/0uWJeSKk9JyL24J69q+POEPtjZNAhl
W015aXN8+CUPwJwddueWlXeJck24/lgof2X1R+oi4sR7SLQnPRlOBDbQl7sXmYAW
OzaHAP09POqDee11VaNpZ3QU39GoJ1dLp22dbPBcKr9V/4KlVqybaD47ORH4HR8c
VoqMJRHV9+iRXkVyGElgnnSpSMBrcmFqiSDj+jAPFROWz2VzxhItkQY4jQHfJvnX
gq4OCSOBHjdJ1lwtmxGa9LkYXf9ibKhq3ns7pEwQhdoKsjCi2+IhF5lyQdzBWMEB
t6B7yGU1IYtPcDYT5KxjryHlxC0q19ehw/9oOTu7NF46CkRTscMAJg8cKA0N1JbY
m56znL4MifntFJ9AzXflHVRTKxBFiJ79SGuwTW4gR/owz8teRhRSSigzQaWRnXbd
Up1QETgHqrhwOq5P5Ty9E5VAGR9pwk92p840l+fBfiNi1FSeQBumDgSxeZN0xJBG
hUmUISS8GvzMX8T00x/e9jTskwxnndDf7BzbAA97LXliuA9yxZ7rBO6cdHWFuz9E
zq+SPA37U9USLD5b8MtWybEZZmKKeBjN5bcz83OQiWnSYfZT6UpPaOWNkByibUOs
8rRKW9Y7TzyOx64gK5JahbOF9MH2ZT85rq1xkxPXimxiXU/B7QO22wi6QGRDkD+s
3YrbERnp18U6QJEObx4dZffL59A0eNUrkShBf+EgNZD8Hl53P/V+sAKAIf28NWfX
K2RheESmNXKgXtajtngHPsR/Rk19t+MWbbkm79S13eLbrMs/y3+aYL25NTEvxOAC
uV0WKS7PS2l7WbitFEjWc1eHxMsF/dOHMY5w+IVTR5AMD9tPjqrZV72MarJ4OSaU
BixHftKvFNdSLwuJpAmH5hg0LGiTDhslGPi7GNGF1YVHLQELsCRh8hUM8yq9tLmH
Mx+gFl6wJG0ryBF5FchFnXcjKA7uxkwv2YLWX0nY1zxFKL3LC82Ex6UGoF5+FTsu
bSQ0TBp+2H00UpYedTzygy8ST1/QULObx4S2YCr4GkPhf3kX4K2ZeP2La/+3NY/x
A1B2SgIVYsXuJE6YSvreJNuiW7Sumtq0///EY4aEjGewxOn0bSwSsff39eHVg0WA
WwA1VjiU+/bYbVmbNchxUgs8COe42iOXzgcaQziWRlncXAHU26/vfqhngVd5iBTt
DhYqBba4qn2SROgeyWsELiIq7C+QehrFpZ08FjxpWT47Ry6AHfYErRojXAgm0s2s
Hs2rd7jyi16P497GZaFOsKxkQQz6Id3Xx4V9QSANc3Dfpj2R4Y4BnpaPuOTJuS6Q
yoBqJ5rjPHqURqms9DbmHkz1dLV5fIpQEPUraBxc4Q3RMxZNb7LJXjFkUAYoENIY
oqoOxBAs10h+/WNgOdk9bS86vHy/b5zvc4rnoBTLgDIYJYNvDzgjEEv0rImbW7zH
mf4lhYIlpJLbzBEqkuj7o7TQoYd1CDdWUSy0LdNcZC+zyaUmduDQ+5bzIy04oOKw
z90wuzjN7+qikLeLXlqjUS/7zJSRkbt4g4QqiBgm8McR12vH81Y99TFNvK31Br71
JUQ+NC7tDP+nuYJ/zWQTs2ooKpxqZYe9oVtDdtwvMOAe7+6cMGoB842t9oQmN9wR
xlCfpaWO5xWyyDHirks/0R1WKFxOG2Rxmo6lOc4FLGGEJNX7U0Xo+2AGJ6TAdyvJ
1WmFINvvXhcyPVdC0EGpKzhlzlrPpHf6nqsbAA37dQK+D4er0HpiIZplQ0WISLzC
cGuAJTsnivWQAtFA4urazWr0kFbi46nOLdeE7qYbAsBxUFtiCk92B4ECikHy0E9W
aOQyLHXuzpVC0pWDpj/yNhb7TN1cm85wxp2FIdtox06HJEEWx3azGlHXJHWUlclD
BkRSg89nsa4OqWxf98skzjw40zhZsPWcbtgOh0P9628zypTjPtRMnqDIza8mapsk
KyZgl0Jy7TDb2aCbfsqy6XLwR93DzI7msNZNLqgE149Mw+A+GSbh7tOWyLvT8TqZ
3QAN4OM85nbYC1Wlx7M2EvueH9UQrnZVmFBwVguuCoVLrFoO7nG0lvTXpTjXflND
1wK1XChbkXfcz0ZTrl0eM5pf9kPqR+tBBHskXEK07aSyACgVMm58cs+RqJqyRN5t
x/sffJz3MbDDOjQ8MHXMdlCEf83FubCW6r65RymgJOWzD3LRn1jzjcPEncFFuV21
U68/ypu+CzyQfwablDK8otLOghRY7stqiszj9lqoT94RH+ZIBhqsUgEHKBa9j6wY
gAEb0dD5g5SkTgw/M4fJnz1O2dAq0QBvhIC8ogPI6QFmEsP2FrOQVZjUHN7idWvR
qbU5GDFcoim9+5gZktECG63ZSSEEGTy4rpQoYuPHA7miDj9L2qmlr+w4lrkMjYkz
NAJ8w637dGFXXPhlay4pU04dYPIy8BAv0bYB1d4OBTQtd89CFTDyLStbAOFmO/b+
dLNcK4TdTcDYT+yiPEgF1DddPNK8lwEBYYPhqRst4/rA6QTYeVoCStQJcXHRV/Gi
j4giYbEHhGDbkms746b1UIxcdXQM56dWTMu/hLvwmA880NLFBq4Gx6uyvDcIxZyO
Q4RvJuwuZEOjP3WzHU+Y6INOHQxWIR2QDBCSX8L/VGRwehDLh1VLNsAJ4gIiepqa
YXyn/pZX8Y4Xx/oMvIZErlP2iMfZbeocLIwMCGTSR7mBmh1TtSLJedcrcB08xRqd
Fb2G0uu32icTjNWqDc8szp5ElLNhd/9MGK78JacmNVsOV7AAC+UZI8w/7Bmvq8ER
PeE5QQrXzSan5EBlRxPe/4xc12ZywooBkVbEn1mUvbEbnceprcCMWJFI3C7yrfrv
vsOJRJv8sC9xJcB8FHmS8z36jMBcr4Qvp8KV3xqAPgdoJFDHLRA/p37FEPXzTbTX
OrKIJhl9pGJUFiD4k1w49ofeDw9CtDlmnbFtQmvRA5RA/DL1vpQbB0wldnk4xMg4
Z13FqsrfWhJYubfPKpwQq47UL7fKM3imHpJrDbV1zEuL4htmLTCN8DP005axhDw8
R+JYUR1PvD2tkg0qQPkSXJKqJGmBpTciF/v1WahiuSVB+CIUrLG0pPgZ86KS0CQO
QCVQKjdWYQj8pAySeF1GvncEp52gTHufZZNXLZq8k2Aj60SmgScnTIEkxxNbfjua
iu97IEFbJSam8uNx23r/aJrmfaUtalPqIcmFlqXizJIanYa9fcDg7noWs/MLua5f
16rJ4/XgALKlGpKY44dwYqoLoPSmcLln+1jpWd3pYqGC2v8WRDx6z/rRNId0xm3Y
Y3QxnFpO3u6bWgcP91lrGGOe3gYnZbbk/5kGrLtPgvBsfpQ8pfEI7k54a7qPAz8a
Ru+U1rGm48H937/XJ5IMX1zcqB59AxpLUuSU8BcBZPegJ7fvvlM+esFfQQP7AJoN
ANWahuGIr8lHFnW4ND+7Nr3vrLXmauN4le5mhjnUlt7tGIOdnYY6pIoaN+fCZI3K
RXBXyyAMKTdN1LfbmrMqy/sBa49arxWHFoDR+FbY1WPsrfnrocfcGa4xBzpWckNM
XgNxdFOYGc5j0543OQHDw1+2iwna+AcZ2HwClJYk/aD0x4KuddoIJdTv9C3jX+lT
hbi5An6UQ/RfyshsU1D7a0jEFzJoXZpoQZBBfOKH9/2qqc2PrzVHRu2eMFndfN0g
bK+Q0W2mTAEJZPGPZz7tOX6KJ+nqXV8YYP33uSsCUypfo+4LQuxgG7VaYVa+KLoz
WBE4UNuSIdgdLiF9tBGWtEK1XOBkBA1Vnns8mVgUrEepntCrzixC6Z8PnjyJ7cfl
eGujIfex3mxA5mZR2XT3sK4siScZYHy+ZwbRPBJXn8iOsfQmd1Fj/uO4o9KHap3H
0tCc53YsoMYRxEJdBLBEuX/2um9a/pNsapfsO3aubO+4FrVUkp6W9Y9pCcC3Q6S7
qNvLUzZ4V0mNO4AxbiiNC/b7iu+dbzEtfPGfNBxZoZMscfazOqUAxzMOnfYs82tD
xppXdY7ddtW9KXAaaLTZD4IYxDbgQiQ5latI5wOSAOZmAfbvQU3HoU4PZU0K4d4v
eRBsWgeSr7qLyFecF1M0VqKVal0fbzDRsX3I49U312O7F0Om+MER9rTV/lxa7Ctq
f8mgmOWIctCAyPwMfIa93Z74X0WKIJKvPK8fsg6Mh8SBOnP/x21jN57H7zGU3Uf0
4hhoLyvvNKtUnWRnW4RxOSHGVBwUFn+wBfr7xXmuCZQwDPe3bFlaOA0vv4JO0COH
Sbdi3SbK5NUuWfuAaYyBTaBQxYnljJ5PV0A6yan3B/H1d8ROaztgV19RuCQBm8FO
LBJ838S/M0qqHzjebzA88EdvhF49R5P2UFoUqX2OAMSPOpUszyScgLEN02Fm639l
FtUiMJpmUpiqbf7cblskGISmv4V8tj/Lx5GCbU9l6eBewH7UkMOxAZ0WKIiDAhzw
ZpifZgM4Cks9+OrdMJKBRATAdy9Ye2NtaGvJL6vsOnzDVnpG2eDEyBA6TAW9hhqr
V12P0+uv/zN1q9sLRE+x/+3ZL4Yjjf4nz4rUamFnTrS2jn7Tf2lSWVMcyREcfxSQ
nroWu6SG68MKvWIEqhX58FG1cjS/oVJE1FKt1PmOiDAbrQdncAinjuSrS9j7t0Ok
LY89LnAl5lWx4RieP0Ij5BdubazPYkK5oLiit15GsvRWaSOTU7n/Lf3MihC7xuLH
3QfYg0A0aC82FbApsG+IbcdVTpFNWeWQhEmOfNTnqjKqZ3K+eOjbgYwwum658/sh
XtFNnpNzujFTPaM5pdYrFunAAjK4iKNGDC0n/ES7IBRIPCvN/p48i17AL8sUYLoV
BzXrHxX2/25rvURj0SIQVdoZr06doqcvW8c4QEEzWyc7QxXal8p9MN6QikzrPwJj
ROzsApnHWkImJD0c9lxAVqQ+e/SJKfYeY6+Y4tT2b6AH5wxo1ZySRvKrH0gyMM1l
qpc+rt4ndjcSmZCIsz4I5ctU+ZXamxZroGYA5vXd+O4x6c7dIOK+CS4ez1IWdgZZ
TRba9LbenAlZKXQTSYa2gy4EHRdZAxLqMcWn8HH51557eQTU1wiJjpI32gWzlSz+
jYKEPaWIA2OiHxJEnaAKkQjk1Kmt0jfse+9R51tSsEmfBbuIy8WW+tzAzzBO7Amy
BZmqXthz/Ul4bGd6di9LV57GUQUj7YlGnI10C94HH6almTSUWQ0IxQ3JhZ+GQtbi
Zlrrfw1K8UEplMEQjDri9Wsb7UdIERLQ0JVHE9gyccOToiVZ4I1mPlEyOgyTImVn
AJenAJzaBkIm+E1LoIBvRs7ayEDz1n1kg3t37Luleghf251XI/GrDspYl9lNCNmq
cdDMGq0JunsJVbB9xBj1hzchU5/ic9gfNTHa8exHFOUlRoBlTcD3tboQE2TZj6tS
kwVulbGxzS995LNYfLJSTD+RD8NMGepLvX9C/Pjj/YujwxhjITqms9KrZofHiprL
xNVZ/mjvQXiisoWFkpP9HfQHuL++P9UguI+DD9FY8aOx5E6QOmmDOxDYo6E5C/9u
D31GhLif3AX76e0D5gqfLsPiDcQNqxSXUBzk1HLbcqoFczsaCoXMVysNoLy7PEVp
kBIEqc7o7COcGjSB9v8pGiNvT7D00yhF8ajiqu12TVkjes0LLWkzg/2XhVpHpU3v
+t5bHXMrIki8l9o96RnsVOaPhu5FFEqfHn0mwTXYvyyv3FoXBHVudjsdthNFBX20
G8QuqOlD6PRnUM/V6rOTcWMzN7J8jyKR0178wxuR5RulJWFihARQ0Dkd02qiSrJK
52qtkFvkWpARekEcDQ7BusQPUonV3/XDPKUcN/V5eXrtH3Gxx/dOtW5ReBE6vO7P
K3ceZRpKe0sL0teNq8uy3JGZ/3NHscEdlGNOFoFPlKn+7HGOIVAUtyp1Bfw+DL+V
tGHYnTpgkp3eOw9jqySaZZ+q4CUB+/rj7fDQeBEnaZZvTeOBf77/LMLd3+4J1MwK
dL4dy4L6PWXs56Dpqi7pqLhau3o67z9KxcZla7FEdvKhPGs/JxZmMIRxBbw6JFPi
ScW0jKoih3XKUST6YhMCJJd6bEPINBQmZ6UTmlVG1OznrtiNM/4MhH03VFaEuUzG
EUs3Ea2TYpZqUJg5kARvZJqvSiOo4/l2FtDzWG2VB2gtUeS+Ctz38i4MbOyO9Pva
ajap8TW2fwaZwmx0P6v204353P5QupfA+e7P2VahPUaIrbBmnWFU0++sWoP05fiE
s/j4ABAzAbF2ZuEDfwtO4lfq+VqFcZJT3+0QgMMCbFq7YJnq+LHcHjV72bfnBSw8
EJNnr7+GacRPH7AsoZC0gQOByNBZ6mugC3T9AfMIF51P3xmGG5W5FyDJz1eJmxy6
/w6jwkO+XwKs6Vooz9t25UdV4x8vLfI0qssAkxCiomjjZQGMZVOh24PKnOAGkZKY
ooSe4giy+TuJ0K48pkST320P1fRao7Rw+d6IGbhVm59xo4NzVDSnSIcc3bYmYhye
/BpxV5Bw95paqoaUGy9WPl50t7pKpmbo0ikq9tz//Z7L/iFSKhNGic0B2JRRzcuk
jYBvHKcven2d+BU8siKVVfgh3fXIA89kVdoab8TSj1I3hbl/1xza/UB/9USFHQir
LCEvFFpKQhFKCOGF+Nu7MjtToLTstv6aozJM/ICZjz4/8FkOk1GbrkqH7D5HZyM1
JMKt7dLVWyobr9WgkGunvDmG4G5sShQ296+XzxD4Mo+kqHm9BjTEZHJ1uFlLUlSB
iqo8pkQCK2a+5Kh0gy91H4G3HWKwcDJ56AGXBE2V+Va5o0clejhygD9eZU5B4T5S
kqBWmudQwv8kfoIk4ctPkS53sqa9oncz3tq2QrJdaOz9kBenIo9HwQQC7gGXPxIx
LHZswu/UvcCqnhn956nE6xIU7obDNXLeVCbwyUF9zwUIWTkYvEnBE6/ynVM1zTa7
sFOY+4Xjzp4slbvWr814UYO4fo+MMujKzJz1QkMJ/+KuTHdFoKC9vBKoEtbI8Oui
omMGAZd+/kDeR6rVTzVnOcShtMl+61A/sEht3GB4TcoTGzO2EzQYJzqpgCrnCnrV
gbyEo6BmjzN+5E9jWg27BH+mTFoP5fC0D1Xjr2fdNl+07jhRdazJD9CvbdRPleYS
Ua1uXa/OG01ufkN22W6gMI6cOkbbvKQ1tYt1UxPhcrlpscpLdXqRvDR0JPE/8bAE
lGUDxeNqYQ9P/zGMxiF13YNWsKCVxrMwKqBNXUVCWAgLTNIaxIB/pP41Zuqc5mHE
SymW838QdZH+XAlw/gSVlV43yTJefscdhUrNUsvdA8yU6avVlTc3O6BuMNUA5Bjp
3RtSwCwInmp8yolu9k/xMOVc8a7uwG0YqTcDJDPyKaob/M6EzeMWTwaKyMl2mtCa
h1NYpZtQW3kCio/1FLdbnmPZJn2fXL0figTagpluyd0JBDsgyI80k9WJbmUBsvOw
WnQOsDWWnaFvkR8WXZaY+4j/8C/sXMqyqrHHOH43n3O8NwsQYWelmA/iXDSbOfKX
MQKfCTGTuxImk3BlGd3zPFkh4OlLVv/YwgI1iR84lJ6a0j5zpK9h62lZ9LqlB6DY
hGV7nNYzoz+QVQi/m4z9iT7WD2yT3DjPjyoTaMZnK7Dfy5aPKCEKf6VbXnqChUFE
VdtyLAfpG8gKj5Sn52/lgpxK3J/qkenbU/rmkXQeLHcjEZmfXNT+dlYHZB32Ssl1
tzOOcGibCzIhEwKwJHZBYcrpoK3oeTrm9gWiRHQ5+HBzrKaG2fD1JMNiPw1+tu31
vRmEPzLY1MMxszNMnOT89L4RIhsofW2sXf/eYwNoi5GTKTty8aVL+WfZVHsx+Mtu
bTXpJY4oiygCyspxJeycz2oV+Se+aJQwHKw9h90djSsGeURa32spqF7+cxKxB2Zp
dhNdf0aLYEStq2sa/D9s11QkJ+dIrGsqJfStLNiL30SSf9WXlktM9jE20k7BLkfz
0soA7GIoHPf6UALlR09RDB3QArjBMUn911j9xlZ7WIZsdB20/FRKHxGKPNKv7T4s
hkMvn+Ig4Y3VgDZObzGIvc0+ZdfQByerCDpcbR/hgPx4j4PRsDhWSv4oamJTkziG
Xd0wUKyBG90tuWHh8Olz8AsBggx9eL8UX7lGq0qI2d5RTqE/IKzbQ6iRtIbgrNO3
YoIhYJdQFEqCy7Nho+yfTDpYT61938JHMbzREgok/kFNhJeEZgTbidz7fXjA6mSA
1rkBbzQXDM0tZEXtpJMVKXtUHrmu/wsMwofRuAyZoVplv3yQTyYG/FpsFE5lVzzz
TiBrdOsP4ZTfvF0PfSnvbvRKaYXAT83SUAjzPa3YCF2mMy7r3ZNTm1qeAVTDPzqC
rK8iPTMXA+G63D4cYKG8xhMehENVYvqVEF/UyBzbiZQGejvv3/cdXruuI7wXxVMA
5q17Zwf2VM067gQYVp1lLv0sH1R9iYZzlzE0TnTHIN47cXo9JINQOYDSuggjxK3F
/l2PICq66M+icfkuKlkErRFai2yjfa1b22y86i+ebb85hJGKV1hsUsshDyT6vG7Q
XhQIW2+uTpqYhX+sHxZe79dLkSYYNC5XHE53KYCipCEXaIqTrY8tZYWcszGLX+qz
sntB8fXNtKyUnH0+sYbwSE2l5zBplGN7g4kbOq2rWFCDOiQ8qoZuGxtpROLwuM4R
RYKZKR6YTI91Wc1eqC+B9Lb+xeKW1H8zBsXeAQsq24VH69IUdE++ohvTBYwJqQY3
0d08QMktjBEQc6NAv+pxtrAGyoAxVXXTsg8Np/Os8fMY2H9LjoyS/XTviTr26uuQ
4GSOuupsL97EjeaoLrrZXynxtwYivQ006iPhGnnqFTTzFgf3a7cJrj2Xdfqo6WCv
5hcRMyRn+ip6x+heYakzg9UTflSFqeTD1K/LsjtSRhAo+p9lDqhXFJqRGITPxM6p
Pcxc6rRkv3Ygj/kYeBRhC3q23ham+bkcDy8586bDKp4NNTZmCLvzXCYlkwSRR4tb
AQwRnAyrAkORN+EhrAE0wNlIyfP5hJ06jDBR63FeNqM3YlBuL2YPLDcr5T/k/p7X
nCPq273ewtMGqFdluZseuWtUdzf3eOhDQGpi3U090/hFG/flLhGZKZWugUmo1MdR
lkZlf1wrsAC/d/tFwxqTUdP3USXnLLlluUzm1hXn6vbe6ita/pwL/xq4yLj4oI2G
YPiWJFylHOIOkXPfVo+kBpP44EVdxm0cMjC0k0wmmxtaC5uNTQeuSmeDhbJxfWbr
mDLh5m2qQhKqmQtKMR7xvGsW4357YLMJDyM0n2UAbysXB5TKdUZXsKDFRStiAQsv
5SNHR3sNLG+L3qUWk7V3/SI5DSimtjcaw9unScgDNbsg+dX27VWIu8yKqlrbtM8l
GENM9hqa5jjPLM0M2ATHBYar+1M4lKdL0kkZER7kJS2dQjK6dAs5puUAY4eGojkD
mRH/6tMuU+l8ls2RGHgA256DEY8TkBITPwhDd2FGTZz7RCEdyf5go+/yxdelPzKE
nBfttcj6eVn/FoGVF+xMVxlyRggK11elExQl35vQ9dYPtc5zqbPl5dx12kBq/cqX
7/h3v2jm0VWJprWQGSVMHvSSTdfnS8HzVxQZAJNF4rUagOrxK6jTXy3dmBK+xvi+
q1t5ucNQ8n7wWMknjQtHdpusUHnQc7kphPGtxwQbIDUWD1hOecs5BBj07lj0gepM
gcji4nZ/+NVOy1+1GXnCFspklYEPrwRPZFEYZEzMF2USSpYGlbEcyq3BjO6p7Jjs
9E7GOCZbtig31ZLl7vqesJ1cCIAM/lXh2oY4yUwKHZgvIjRJK6FYgG8nsSaHsZ+n
IOObOuaTKdQ+ITES5aAAyCfdiThyozgVQSOVEhVNp7mSzi3QIbZIcdfgfVRtIqzR
OcPAaKV0tbWbmhObO8S5S0Fh0DJz9VZwP3vfrFQJMMhH5eWHzl27Zvs1pxZgOZpf
I/4g6s6dhZoIcMa3wlCf/Lh8wouf3H4ZrpQEk6d78neTJcOzvog8LCFW4ar3oTgL
Ql0tRQ8EmZq5B3HdnCGpFztZHIF7ExGPxzD3d/oW4gZYzs1NGWp9i0AVJkZ3ZB/5
gIJ3bXVs5jS4x5eYQDZBuUynPIh33wo/MwxX0YW0mV2P8blhS58QtZE7UGZYDEc/
+34q8nP8WgiF8r/pi0zN89/dQZfN1smxUdXB25eKV7f7wVOyVDzP/qrNr32hhi6x
71bRLAN/bflIpPgHhrQpnTnk5Xr7rniWUKIeOVOGFEszui15OFdcrg99ALSSjrvP
WE/UxDvhmTbX+u3BDgmkZfD4UKoNPTkJYCRljSCkZHl3Aa8V1zv63Mctqgq2C29f
sZ93ATlHFbHIEOFdT+xitc/oKfoC1neKm9/8ndDGmcttWyrVDPTjxG/NTwZQerZA
QqjspP3Pa0Ky7jxcjxrMOZ6n/XwnNycqUfl6qYdFb8YhkxL058rJtmRkLhAbLw7r
4YArclVF99eULezOIvUQMyQPkit0UuBynwmoypwtOflAJyKDSTA+6dGm6PnMJPPL
QbaxE7cbgG6HpGT4jxyCGRMM4kWoz2wWVLv4QEPB49WrrhYx9lQvxZelZCets2io
4ou4j0ljB3tnC00iU3zwQbI+O8WPkwTHD2X9xE/8ldZgc9cASWcoBeo7nTXUOERK
maeUrS8E7UJ62bew5NBYrALacfOoprTj8702IA+KbebE8mliYHcJN3SyELExvnhw
5yscaDqqeuL6SSvSEGLSXvBsGCcEshSmnU9JWF80x+Y+Nuf5hQvmqkwS3VhDZCMA
4LQauojZq9mkEvcKz8JAAVFMLv/I6Kf6Y9xa1QXIZRoLDX/6MQ3+y2aayxSjueJ1
LDsRTjE4ezxF/gmDKFKame+/cbD0B0OBMfYWbtdU4b/HJsnn0lITJrMrns5zbpC9
a2KTrYuxBkqBIKsGXJs1D8r3NYoQtqurrvalE4SBV0VA/IxBqAPV8i/JXZZC0Epe
nlojmTefBWR78JGqdATpVT/GqBIKnQLR0Z12gJptmppp0FE+eJGRrKBs0ttuZ1n5
KGUKMZbMOe0nHK4CISqXRF3RRFbmpJ/Xw/99j1KzlNcTZAC5YK8EMbmPtuyWctmV
R0aM7dUdwubgnmS1VK3L2cvkqoQCGWZXJ9UVApkgkP4ZsYr3vJUpbovKvLHkF2ui
uC3g/fzmEfGyKBTdSDYJOvMF13im7ESKgmWgrxOJwgs2nT/vKS/iXEnBAqfbJfid
BjNIASLZxi8FcZFTgR/JHKHDkn4HtKO7blchA7JC9NiQ65MIjV1Z+zAIkI65Zhol
eDdDI55tvY7JcbIFuICcVjozmIpj602AAI7U2LIYrhuViM7m1JvAV9Zdvw+cLDcL
+cuJjlTxGzC8rCm3U6YT9HgvUKQMjhjvXCVjoPy4PaIX/Diti2/EOr5uOvxt2C+8
lNOrA6LD43pH3SSRQNsTjQWPocsoq3F1/thy+I6jBs0hZ0lS6wC+kplh33w45dhB
+0eyQvQNzlbX0m+JGz+wfotJZPSUxBYJAVxg0Ij6mydxoRLZ+f4sTqoTbdulsHk0
oAZ4Imgl97Ol40M31xQ7wL5Q6m3JWrj8gziR9bEV9WVog4nfM2gTLFhVz5XtxvP+
lg3F99IYXO029shS5bNyJso6J3qy/Zr8MBo77s91qPKrN00wMSA11EzwzJty8JGi
jYrLw6X3RTzcpTbTgqVURS5Gkceb17OZBT9+TPS+S2zjqU+TASPWWqswA+bgc6l3
HHnMA0oFvkkiiOZ/Ccz7z/u1MMip+LfniWY2HsIH7Ac2Z3FgaYI1k7+2Tt9gjEkh
Hw+G2oE0nijpWIUP34jshGV88PCb+vsgDzU4Zv+ydTRiNOaCtzTy8nSR/1xi97E1
yW6TqvbS33rTbegniqHiwAF+MB9D1FXQ05ohTZam3jbp49KseBgA6swAEWYDpxWz
GwSalAu0Mo11rvLfTWvkndLD+Kdky7Fk6BcKDvAe014OTf9Vdn50/vFS5qVEa9rc
IaOehSk6Oc5SLihBqjNmvHnTyBH4lVishVQe/slK/kgWpq1y692e1mEFpZT1tZdW
bkH1EG9Myj7KX+LFVCDgwF8YB0KbcIPTniJi3jZOzbZnImwIka39fLuJUmhKvbV1
yEHFCaJ3WvRS5cbq1TJ4jHO8WM1VDYn2qvmj3M/N+LWJySC3nDYGcrS0sYbkGvWT
gIVedKTY0qrmIcZTRTtbRMt7dXMdsgMTYFMmXWf599tP+VtpeFbphegBFFRMtS4B
TiMmJkq024KKiiPzpcChi8agc0QlIZB5B7SXRZOolGycXpOUCmIfZB9KHMmwOuXq
y+25j6/m3TbAWdeDaMeYE9wAm7yPmmU2KqfGeK2gRY8d+K9EMyoQlq/2InWkx67z
k6F1qy+g578Q0ZG0ZShsWsvk4o2SUw/N1NXcpZ2KwPD6JaoET3FWUVSVnMAgY9c6
NrUMqAdjidVIc2mdXslxWaQcNUX6vgbMwYXKAJqtv7+iQ6/TgNiC+9AbjaeK9suZ
IotEDVOodHrD6QsQERsxdAShAsO0RplhIm44rpc6llbH4rRFAGwy3+IIJ3wBQ49+
1Klg3sUB7f6QOcculRKEJL+aplpKaJhX56WwwfRSqBdl7wdx4DJK2B0XMoL+oaMZ
3Z1XkfclZPN366P5HUplFWHsRptaQMflDU6VNT9WnItZIInGvOo+xezzx0V/5CQF
70GwgXrfo6wD8C/Htm0UmcMQ6e/uNvMT19EMzftLh+ENQ/2rz13jCcijOVuI/pb0
1PdnL56e+7zXpS/Uc6NW8gFYW/U9n/Y2A31xGNZxh6Mf1ceYRswCUiI4ZmE/rr6K
EOAT1/XyHvKGAYy1/PGogMprpxahFu2rmgNH+pt5K9vh0cwPu9UZ9oZrVOp2xQpD
caiMIJjDaogpD5It0PXAL5RLiyo4U9nEdzlcjbzBd+SB29Z+CgctejSLAsxsc+ID
D6Pqpx11hothUXlaXLcheR46XX4xASar+7XQKQwlyuLTlPDHQKkOVmo5ALKbWGB2
cMosrwc2kaowv2zJbrkuEcQAAW+QT1GnoA+GqsvN5R5cHhQXVghB0XJJYJO4NFVs
7t8Wfd2WOeRjOHQ4Fe0ToEN2n3xqWocJrQkzdgo0sZnEouuNelluunS1/KOtPdoB
tjnUnIvTq4c7xCEQRV8bR9yIkWZkZ7vsw8KJ0TyqwpytNtKvRCFCa38al2YKr3iG
dPn0pA4u6EOuNOvfXQRHWF8ewpIyB4UFN74YYVlmi3y7Xrx/k1ef77v8Bo341gjE
Pz/smtVWrULGLt9UBDLHyoPqzI4An3uRMzw8PMfyIv/hSeu0qD5ROZv3L49Emvzp
XM29KcdK8ykQ1zYogXMaQhsDsk9miV9zAEmqLha8k1/a/6bX/h6/HfVN0FTvDy1E
M0uw6JiXQhxJaR/GUdruOLmNpe9QyEp02mxpfVMjP374yZhKL0pUv7A9c1RyQBH3
0xwF+lyVJ3RNPI0sCb7BHf1DeEz/BMWHPh8qP4gNBb0oQXmU2UKsRbqoKTlPgquj
ebO0eYxYNeO3cXqk8wspO7Q0nVQYNqsEKdCwNag3/Qc+4R5W5W7aKP2JuiE5n7E8
nlxOrVGRMU24J3iwtUWe3Ng2kB8Fp5WrJ+ZebqtItgFGYtrCmZgYDxLkk91eQyHW
h//7bcW2RnOon6RcwLL1C4AuufFtwJYqg8xeSpil53aSZNGmxtY9n+upozAlChwH
xqGponUApUg7dBiYSX50CzIz4+JNf0IQSYPI7XIFllY3R/ovWoX5Luyf5PnUI88g
zFvzTHN6o3p6aEdbzLA+MkRNUb1WOZDixPbJg0shKidLVR2lb9fk8wByKOTxLi6G
dsQILgZODFMF8jXyQViAk94sSPM3XNRe67nwzcR8iomwAZlzH5ZATL7tPvN+8f3T
opI/MosigNH4nUxZD21qij5XfxKDbojuTVHfQjjeARGyttRyLKTDY9aE1GUT/6D3
EJzZaTO8LjxrnuXMKTLnJ82wfROg4ysBbPa9xTwc24PLC/D2RucsWMREEJrX/LI5
q5D07JBLv8Mh17AtPEPCrTPCSAmoTq+kKhrMB6A0BNykj2ULwJhoW0dhmzNtp0dA
JT3DS9Mrhn4bsS79dqBGmfTayrH0ntYquvIFhG5ruXaLmmWJTl69VSlQAGieI+R8
rJxewvaElURloALGRmBXO86mKb+Dui0VA7Vx8qlNfgqosgboyH2h+1Td6C/sEmhi
U96MIOTMWxfN0xx5x6BReUDMoxZj795Rv4QsKbysVARVVCF3xJUYcEfbgfXOIMoZ
8z1kfYXPVBLctRq5eyydDHdbynyKvsr1vw87OYI3f0G0aC/KT2ndBZWVCxzFOnhf
04pHdsVHE1WVmstRBE+etO2nrZIuywZu7ng8CVtRFnC7fCYloermAA536qRIZf2n
84QAwz81uqBSTMd2ntQqmdsyzpNV+cWWiTDEMxdEx0wdMukMaFzmvc1WhLdEM/Tj
DdH6cWYcICbI/e7xEZuG4HQJIY0a+4jSh9UF6Ec2H/59KqoLMLzJHNPSfDcGkH4Q
rC+Hx+4ZBVjdmgrWhSfzV+3DffIHPr/mY0bKaouOu8EJznbfLxfs1qbTnWrLf8Az
CoO91PDDmAtSI5CjsX+7nGgUhrWfEdkN+24ML61avn5wlbN/Mmp6yCY4IflPQ7Ww
xeEEa5XSxflKJfXXxKiWvMH45tE2QUfs4cb1VIgZKyi59UaG0SbJyTzV7FQykfn/
wiPUEgBrOi1jjkhYtysZZmYGxc8VnFMla5LTzi9DZaZZQY8UeMycSkBSBXTbT9Wl
D3U/ODALEY8AjaQQh9yAmcyT+yF76DYyUrybX/1ElFV2astjUASzrcQmx2Z6NQoN
L456KwP3dfNTAZZjvbbKl8N+T+HlSBOtqrgo51TvRusw8bBrBWUnLKhswqOrqVMp
Ivnlvt/WKD5M0f155sZHBdZNVfxL05tDf4GTwsxRox9JKneijfnJHVyCZ1anTA04
WxUjuG65W22ocpBhajx6p5yFJkjL36DY0O64gCF+LgUXz43Ue/QX4ye7hSaZhoNS
CcrdOMeTJCAzxoz6ZGWFNqZRvyDDNCot1P8oOLvxelIf+DCpK62lNl2K8/qLnq2C
1Svwj0mynAQrNEv2sR8Qz4iMyqhiV2KWTxOMleVhWaV2uTZcS0c7tTjkr5YXh2m9
4QiVVxHSKcZ8RVDD9m4JgUqzDo74quy+MY6UVJYBWWKKrkG641Gn1p9gBR9Np62k
XjHwPMuHTrG2WOcL1H2C7FNFtd2DXe+Qgz9G+nsR+b9eXjJZd0pg4s550LU6aLFt
5npflMQp3p7vB49O/xGErznHP4MNT60LCemgUrQqBIBQlPsMuhRPFkQgU7CW3M8L
haUyzKjX4LKIsZX8J8k0Z5m1BtCa52aXP6a1hY2GVs4XzllzbMUGA2mdFWjAUeZh
/g36iVC/bUmXwrhg9nSY8hevXB8f7AOeqRTB6dSCcNkFkNYAsdh+lID1nd0LRlaV
/8HSbeSunbBgFaeQboC5dPAWG20uVT7+Q9z5ZxdPJmAgcpFsRabKzXPE8+Ta5yBc
pmyXEqrNL0vEPeRmnuZMJTV9wLSgQwWN2TsZGH8RPR24z5X5MuLlp3DoJEmtPs+6
jdncqaDCHNcsr3TWhYLttM7+o4vSs7amzXOYM++ISv8jAeJAHuE7TE768jvGsd3t
bDTcuLlfmvWvwDscg6LAIk3f4iSWifrZLw55xgGtWcCqmbKuUw2uH9SbckHJaz1M
qQn1uIswxsL9V/hNp+axIeb3rOPfdQ3WQXlUFqzmquQw7Raoh0a+3B7Mpg0fGwCt
raXzcNIsT9cE2dTZ4hm0RJndy9R0tGRI4e9SJ/VQHHPkWkwR/dmSZrBWtC85GfPJ
NvjW0uU6urJVflkC988P/1lHi1IAhEMl1Jd5ejtIjy41nqf6pqy36wbUmTWuFIy9
jUISzpNbqe7yIVR2OUkoFSr7/lAYuYaNh9KNJ8qL/t7mseREffg7GC5ndtVBxvt7
fdUG+SJ7vheSMNZLwESIdOApfW2CpV+pj63kcFPH5YCtrDRjfD4bIWwXXbG6pbOT
WL84iYdOX9Up3PfU2nevTVmgh4oGuGw0KfYOCcKJK7WaQhY5xyonnRnDO4vrPgKd
POq5iUeon8MJ4xLFGx8uBTtVIPWeYG1Z1ZMrrS+dZGWvkpdV1DlIWIomWNV8hpk5
E6lPwjhjgbUyXLMT5q3Ye95Dtl0q749nsBFh/GoT+SyGsEjhzlr7gpj4ch/IBvOX
GHZXsOeGIwjQ4vAGZYh75D5XTavxhBrP6M8nGJpelPqry4X9LEkrzWuZ9tlynldD
BioUtHjI9c0jSgz3Q4S6tLAWZQdGjAbmp12ps2k5bE1nIuXNTk4NIdPQtHgUoROi
i9ol2Xpl4x99E/IQgXmgStkQgSOZDJvrX8s4SunBF/qi0pPVDtRGScXMN7szDMVL
L/sm78Fm3x+4Glti1rSNG3oYaUts4xDVbKqK1KFTSECJVaRZ5N+auVLrSnL10/A3
52zswRaOpJDknQM1xJatDMJT9BCaQKMkfm3UfO3uwdYLD9LnEtfCsVxcUWJUJPcu
AsyFFNTH7Z+bDNSbcwAm806utGNonCqyaTiWp1jRmV9Gr7Jv294MfYOYYR327I2Z
h5364GtMwtp0iRan2gnOgVPqgE1dX4lzcMwAc4eZJjcWkTqwXr6vrY27jf6G57fj
6GgdjXywwpXd6sN7jNH/P9jofEu5osx3UEeRmZXmjhcd6ETMxEVRnISE/oPEumbR
wbfr6ngM1rMkWL4IWrsNeMEEeXNnV2Hn/SwzpNDLLOt2T3WMPQeNwpOiWPxBl4Ie
sQuigvfKVX1HlMHOhXmv5GThCfwbVJq65Cksdsif/58kM/E43qbpF45jfFMQOjHd
i8jzAan88obhbLaZVdiy/juSfdrMgLZrRaNJW50DmauDFLYfISTyCAPVTW79a7Lc
56h981QZisFJQYhVZ+uewBisjNDOv8z2VhhhHMW8FSwwLoLYl/qTRdzaMpopmEau
sTm0N1jXoyg4fhdUpaX4Jx275PxRTmXFAm/0Qb3jihZ9HvIe4wm3rTA0qnNYACyK
EMwD3fPo2JkuHUUbNqqa6VZVDTgs+K6jtRKWN1Kp/sFPk1tfSjxtUhdkiecDD9oD
TvpyxHiua1nuGD4W7r/Gjiqe8Rkr5GLR+CjiEOBWETNeaPoOrGsLc9jxzWuaCKSN
Sz5sEuW5iJHln/Fl2JWPwneImG79etPsh7Tkjt3cEl9u/YGnDp4f5U95kcFvvz8M
KIGjNQGxHm2/PI/1Uc3zP7olLhMHBw/NYFtzjO59ArTeUUUh8qI4sy9KvN42niT4
mESy/mAHLtMQJKOwHGfWylDxPFyJ+Cbe0GlCQ/LGJleB7IucxaaFvtyxUJp3czL4
xIs/Y02pI3S4YzKnSBoNZ5CsDLyIbBA7JRsCpHLd0Uj41yw9YdcNqZdrOV1pTXZj
mDgmsLgbXYLgAQ1JJQoHUI8k7g8j6+kdoXKbFtArO4riuZrpSke10WMob5a+UwlH
C/sCBGZVB76YXzstpBs0hMMx7WlHQgAjXnBUtSMRj/v/xCOKOBDGrbPnZ8PWlYH3
XUs9wEC/bB19wPRw1RV5nkraI97FeUCameZBwHmp2KALlS9hympIQZr7H+7F2k9V
ll3yhYGbR22m5ONWfLBMO580iKBynOLbjjroDuqOOBT5cmczhNu83SH+w0v1tc1o
yp3xUGvFZUx5A37TNon8yBDVd/7uoiVWs8aE7X+4Fn521k9kZtQXnb+jEUgNMV2N
d8RrQKW/zd4Hcx9Hr92SAcT6lllgBoYqmhZzy1QknfUNjx4sbWHzWriZ7ooAhPuw
FI3WnsxdZlhLLbpiz0s2AC1k7jlB1ZB2UOSlhX0RaIeQvVbBvkr/Ytf//ZdPVp7O
U/Gh4mcGp3Pnr6tnfXfohKe2bxTffOYJdUecT8hyzZsM32jRlb0qwut453UuTsxA
U+NNAkD/K+TBotaOV938W2hAb3fAU02RxIo7u5GLAo9KmVZuJnUFtkmdfNKfrHir
d9BWXeQg6sJsr5S4dIA2cJdV0BRVpD9G72mRLrOrhnOT8XVWIAWK6T0hEsuuIPym
kyAuwdqaMBVDYCfrBztmk2w+2KmQVe1hWevYZ/Jg+Y1oJqPQpKXH14cP7Va8XHot
qugEVKAujW8qiWuuHidZ7aQa9A3IwoObcB2mL16nUKNFcEz1cIZhGDyLSPX78qEO
hZBKCDneYoccDvIaIvaWE8vU3+1onvHPGt7vUXUA3/wkPRKoloCDi/zJEH3/f9g8
2N2Y0Hkr/ceTcHG0X7DUtxeedO6idz1rlnDzrv/Sk4jxrsts80dJaf4MlzT9P81c
rtDVab55H/H1i6tpxBGaZK10oTTyiD6GaA1bJlEkmFLam6ijxgTW2TPFYrEe0uhF
llJUP8nq+6DlRFeSv2xEb8GU4S8D7u3o+EQPTmHdUhGX64aSudnQxpeIUDb1O9ep
gi4h1WTu5WViIYdIWO/OlP32f+KgBUT07jyFMny8KxHaEgjAKjMYnElm1aCb9b/z
EZK2VqiYRWoLSD9KPoAjdaflWLXzU80KpYFHsHlJvZKgm2ZNIa8/hxqY+KDLusaA
2TdKdD3nu/iP+DGV71uCFvQu7DQNIbY7K8BZ5TsjJcxqAlg/ThBntypxJ0OKQpl7
IwKCAywrWT3xKeEIr4oovA81Etro20b0CRDm1S5LnoetsbVHcL+82K12wRQw0KPK
AxqCXR/bh7slYvwjo+30gwN/dPUTKrnou9PHpdFxMfaS2eOUFghYdxNiKfQuNWBf
PrbgYFJXJN8VST/NJ49Mc7szQZnP/AGlp0PiNlqMR+XvRAzmDw+yxfaj9HcgwRmG
7hoP8LetctikS/UrBE2fJNhR1T6RojQulcbETwSu1XsVjBXsuEJlwN5Z+AiLc0Jg
Np/lACJs7vwdPTL1QHFpZGsHUmph2VjZ5B1MjnhrEsx+tFDL8I0rpKyIi8+WjcXZ
X74NWiCuV6aoqhEQttud3j8NtCmSz9V9FVlmPbDaNnQkdgXQD5W1Axxiikw6j++q
QSvdSDZRzXyy5tAvYpsr3mqvOSktrmFyoy9knRiY5W7cCWOf7M5fhf8I+icmnBGZ
Ag2XElzSXT+uxukS9XjGHgjcQSbeX5wyRuxJOOllwPgYT/Tji6S1Rw09yg0dl92j
NsUcr3lrkua2Fq3+AMfywoednP1sFrguG3J5hN8qIRDGGPriGqQBEwmp6rtuudul
pfoeE736v+yVrdZLpv1vGYY9dp2mRsWSugT9NBfrIenRYce3Xn3jGLSa41oXh0c4
C8w4CNfOfm/xGqrB+heanRSnI0CXxyOYIh7IReMIwR1SV9fGk+qImg8nGOoGB1rL
748sZMfwMcp+yAHhbLnrKodRr/mGGyIijQ+zuYNVACntwNhx90CPSCZ2k6GuaGTz
e5nOxhMqgP16L6t2bWAFOD7ufs6JgF/amhezXvHPR95JEAV8mpB1/6AGE4S6F63L
nOiBSNaCizO8UjVAjGUOHQh81QKBEfcshPjr2NU8ERlByxgUX4euzOtZj/Xgpa97
AOTCfA+Q2s3GczXi9DHRKcu6XHIezFAJeZ4KG2sLfLs5IQn3cCMGEbPuHrE+IDPA
dV716oruQc29IyOeOEmYljkyEkbe6DVvCge+n1Ps4DjLJsz5U1a83EBvW+QjZPyl
OTlhvuXsK/1uMxJZmuqHBOR0sY9W5PiZAfmOihJXlvY0kOPX/fSl/jPrV+KhX5lj
0fM6KbqHPBFMFmPmMseoIagcDNOX+F6AvKFCuSiXTe/t5oAiNbHptV4avgR8oUZ6
t1MOoDPr1wHbIZKETISCpN8aJERoyS0s6Rt28fS/GK1M1kIRCIQl9tlOTfo+G6KP
Hl1CCLY5mebalGO7C/eAkuIxj1rUJ2QNrajKqbRqxR4IqBzlcKAYBlAIMyK/FwUh
56TuRSBoEzoi33yVlPaly4l41H1Ymy1vFYtvaysnhfc6T8ALJxV6xBr3mLryHpJk
9v30y6HSePkZ3D3x/V8J+oc2KrlbF6U8XNYKDXuAaBrnGvAWVkK8D+eJ2pSPCNoi
ob5z0TfkR3MnnuCQ8BnAkBAORf8FgcR1Jh1WYIDjnqFZWMItoeYC4KC6/Zac9xwM
rE2iRSLSWD62X6JoD8lyrP4VyW+6lJ4obgKb1GAUegULKiuRZ9BAQ0RnInhBgAst
NvyGpBasOqBbihIgwtUo2PaFHXunU7t2ldfFkOnj0FufFqiOmgTBirL0DPm2p6K8
ON2s/quJtan2Z3iym0dIr8VVjQ88SuQduCeokt6J1/LQEoLFvOMU5DqRs8nVEC9L
m/NHrdKRzJUQgGYtrgbD7KXOhZY92lkQ08kEoJINup2VktJAUiNBEaiYFPw0qJI2
9L1xbZaOTlp/poGC3hyfgQyu9ZF9jxtJcogj+b3zqyVp2s/nivYbFkQVPS8JUaKP
XdCqhMHKHxtxx5+PjXxGllfIfJWA0baRe3fFuRm+E0MjlAraVNU6jhB8mkUSLNZ7
pGyzY14JMqlzQP7y80XoilpeqXx0nhGvcnFa7b+3TOsBsTdX5EHpCN0WCkRJu7C/
LtZYPk/64Cp1M/Oop/Ver3SLX0gia7rEhJhBv5cDatTzx1rmBrkfbQlR3nUucTmj
zN1aCG8sIjdB0lan7T/5cwwnGYp03yxwxvFkCktEfu+LuSyOo9UxtEZIgrU28GH5
7g9VUZIhctygmU8vBlunBhsqKk37/J2Pr01rQsn1waI3JWv5IIf2JanHmjGyMRXE
4KXC0+nR6l7qkFvXEXrcHZi+6eqrwfB64WS8Iy0Q01MMgPXo6oDHmPLx7DpUwJ7z
e/FlP4YeIrHLV+7kXfwaz5GyxQViG7JILnoOB9N4fy24aj3toJv6tH0v06LP8AkJ
slCO2VxgQqKLDGVCfXeO7NzBOSwvscqjO5SWpoqGTuZlzRBRHp4fM4wF4LQMqKMY
Jjjn1iHA6A2WIBG0DlQdTGjvYzhWd20w/an4hF0NmNvKDPLcLuyQpKw6iYc0/vM9
EujRu6iH2MDZafuPnT1RbcTJL8K1aBC/cxFPcQCj6qTUdBSMnA+pxFDJX11qUDdr
KMwkaNNn4F+tQ/MJRtnRRGT0694o6hvGWlyXWvI1aW1KWkCcKU5N84vQSWJA4x9c
lrRzIiqhxH8yAAKK+mXLdYU9McaFp7dUdlwtx0qK2JHk7NxYewXqNYwvQ7gEGfc9
S+JxMocO0PfK2+2+Ap9L2irZPhGgiP++L5r6cJYfGbiScYMqbSa2oYnIKdc2amc9
UD4lJzPQb9NdXAO7lg7xToCZ2oA84+Vt0Qf+Hql+TXpRTC7Y8ksHLtdgwFVr2iSs
811NWT8ZknkeDjtDsU+3h/TkDPRvDjQVOIhBx6R/JHklxfDTuBBbIs2HTunX0Sux
yVT9YzUvoLwJvqvJ/VQOdcy5Tu5CjCxw6DyDlHe+NTjArt7c+AZc4NSbCcytdlZv
hAg+xCXySIapX5i0N+klsWnuHcyOAzkR2To55UHI+mucI57v7pboUKB/XE1Z8lFt
UkaHtOZFHUPk4PhZ2nkPeeWKj/kdqn2SuFypDjNsDSX7ppHoLJ5siasdQL8wrU+w
NRyIx6KToSiOw1qv6UWeJBhOG8VX+esB62JQVdKrizu6s8Fh0IMl4eDQQWx/DPom
2tDXaCCBKIIggnlPSL+gvJ3wuV76NQ5Y7VNgXTKF5CkGV+wUqjFbE02FMy89PtU1
dYOkuvGN2wOvTfzSoMcEBhtmYm7r4ZWawd3bMzzC/TBGuSBN8HMOfPK6PixTMjvc
06Sf3pfgSVWb47eceInwGqo2ciSLWmBCxpNktuLLd/4tTBxHHh7y3lHpfhXlPJ0z
lRUHKXf9VPAWZP1JwNvfLFIXHZwAmH2cojZzH84UW3G0UWEGAtFaELsEI2/lg7vR
XUnh6MPrsuv3uZ+kCSQshV4/KYuvPJj80gUEj5SXhfUNSsU23t4AxchhtJY0xjVA
2/P1dO/iPgGn2YyzLWxZHh8lpPmkkd4e0kAjKZ7PU0PLaN+pkjdnAlp5tax2yaNa
hnda+/7XnBx6izHXScQkNRT+PCFqcKD2ndnir0i+VCJh+ug9jtvYIQQodrFzep6K
zO1x3pmr7kpKynO+5p0nTcJeLGI+lfSZyfsqQttRFUGnOcIgUuiKliRt8OrwPosn
q5+tBbRoeo0nriwKCZRp0fE+1SCB2lcq1HH3i5Q637GJ2DQIpbkK4ao7IPbXjs9U
ScwADZf10KA/4X+WovkLR1CmkRQDXOascv83KjMpDG5S3nOL/L2Th2SJd/OsXb73
8spRHR/x4MrjvFOLr+NsEiXdDC8CJvWN5va7ojbwuKM6EXOPpk4uDcy5a5QEIttd
+z86J0sSZAs5DHc+XBcm+0NGFdd3vWGEu9Ym4vn8al+fvmLypF5CK99MUDLZw78d
a/qjGSPMxhYRSLxk4P98G0gY7UiqegXPBVg4x5yHD3/oVCVu7S42u9YLEXMXPI+8
iWAczGaKR7E5UFKp0aXwjBH4v5UxVj1JEThGyJlDWZb9rBJV4WGwjFnen7uiSMOE
WANH2Pj3U1pU4Z7y6A0AV816Mh2kYRsIjtDwgW2UXxQxtPS+4FHFuZGRPz6w6qTN
LIoiGx5SoWdz7nRW0HuldhG4+HCof36C6I29TFnq29dHiSD7YsxT1LMm64Ac6+QK
7EuchF83gsmjSHjTjtK62yg02QQYdQsqeb5lHrtRdqs5RgTQFApB0wucUq50P3Xc
PTyU/ikRipuYecdFbIx17Q2Bll4L1+vK9XKSpr2/5H0ux+Dp0/eYf0+fz2R/9MvQ
uz/yxELbCdxWt76IVcjKb4qP4uedxoL7WaGHeZxgxAavt1aAqe5nMITdHcincgU1
3rwEioyRPCBgjn0GkcQuM80b8kCzmn8p21yMV+psglYb2q38vlUrPI+l1FMjMSe1
09zYvOVo/1pQZmgzwfZNPHoyrvB7NCSg+Wsqs6PWTkbOYnwgFdQ9U9/m4gNlmWg9
A6KQskkJ7R6WpN5rs0Jnu1k4B2MLKnvT6jWjJfZ2CT73tCTv1YXtfOaXvdCdZP+Y
H0a9rW/Y+FNOeKy07akGCWrwbCyqUhqam6DHdg9ncAlp9gnjI/zqXwkxbxV797BF
0nJ5Rhn7io2+xZpjxVZ0bEtHP9GTQpWPX7+fXATNF5pBTuxJqEyHzMMbM5IBI2l/
3UxcMsFczKddlZcKLGRRw2ouoOEhis/OCG8xh896ATOEl2uTQH6fiyi8islZrZHT
ERrnm0YmA7FVBgr09otg8tVU0ThVZCa687nr8L+JC2/gXjC8Ko68KdwQ6C8EPYYF
F20cUjf3HVv7vN7L8l+ZtyFlA1NuSDfBG0f8l6bZ5dJzOMYpHJTsUIuzw/839tks
zIO8ZnB//EOrdnb2KVHwKXf//CiVAJMEV+I1Hrl4RLFPLEuDb3wCK7ie/wAYZVZN
GQugNTQlyIUzHx3yl3UaXCDu7yNpsxhuE2oLHT8X7YkjzxP4xuHU56fGudXV94Wn
xtdIucS217AXbvuwlF6yKcQaqSl8X9tVMZMCXRw6qM3D3v8RDJMgL1mNqtOy+4oM
24MDCU/fcZ2D08pM34rTHVT3RmmNJczmaANzVGYqVkV6cpoLOL8blP6Gp3/4Br/a
cexJNHfw6aMfHmogPIoRR4RLVewC/vpF8zoCvzZVUz2usv/qmX0SYFE7kltup40v
5ZNGV5WmVZqdbKVLbpQFyhFf3x3bo3M2bbEc2sAzQWulhegr8Y9/oWrdiPQFhy7r
0T4NSvAhPPbnqqQi3ArdfCG8fTjamZg62yQy2aoBTYM6EaYOw5dAVNPN/V+B5O5x
LeeYztjr/aOL2beRKahvFzU7iw1vd8AJyK0QV7L2FpnktmtTiSRCh8eNjsfeQOPu
UAzK9I7pqDmT+yUgcjyOod/bMuW2NGCwZSfAl1q6Gkn3P8HJKinxdONUsltLq92O
xGA+tYxjMrnSqeNhKWf7g7ZshqW19/VNuweKplA+bNMK50RaZ+1FTAwH+kd1ONhx
y2Wnl4sWshwf4J08bM3Bwux53r6nsjQ5xSfgl2pVKLdqOcVwjzqKW1EhO9ZJSya/
tk9PSrWlXa0bonCRm/huu1YK1BoAAiV2BPUpEvoQKzI85AAzWVMMenQ8VvDxxdyE
KDPzTjzJXG8cfqe5U3wtqx+YYOfor8mJQUQvW4CeTth+6FitLv2riXJ9VqmT8oVq
ukCX9S0GCrHZTPsEqv7XHOXTngo/6SwXmhk/qdp9xyUakBY1bjRpFzU+j1bd+bkZ
YOFaQb36USAxseJZd1dP51VmDFnWu1CLJxhtUFfcqYwxBuj9qA4EgMSNBIGOWh3L
GdcLZ00WIQ//g3LBKpPERIs3RKmbOMxtxHY+iXxHrvBQo51vDBvJRxXckdko5azY
KU3z6MJnG3U7493UTnr75wiRY1XWEoJQzMVu9tv+8Cy68YigU95Ryee4mGYyZqPN
d4378YKrBvy7xcv5Ddps/D9KgcZH9CuJe1QzYS5hmUakoRl+SqRwTaeAHd9V+kQu
bz+Eg7M4bPryqkmxT3evMafAtj3BNi4AmpCRZES2Y+sNMYoMlnASscYFmRjtWtfl
RMbUd7a2GlgnpY8b2R0rq7Gx9GmstiSNiekY56oC6c9GMDreqBMKpoqTpfkkP8gW
/pg72xS8HlbWbPt3oRtxHIbgJ3T9XOoK36rq5JfJCe1bmoYVu0OVQ18F5mGLPrvf
OYU7sZtu0PnBnEiuJkvA79H1m9OZ0cf+hSj6+/xK1Es38TCN4Z37SbbSJIxSkmO0
D6ii1yZ45EkEm9WbO5UQdD2aP5A9wOKhcPiftyubeSgVdpRWTQhsXE6hs0WnEBaq
iVPFkazBOjl3+ZwIZtpb70DkzqO1Y5v+cdYZ67NC4DC7qJdKz0N7ce6wuXMOt+YW
0WU2EnxxPufnYwznAVWs7Wpfl8ZnaF4UNLe2XKqWn8+Qz7JKmuq+IfVEoUN+lQAY
/t5NqziFezEz2Nq3XDkY6+4hYKdkgFrmr/1B+LyLflIk61b+aAmSjTmd4TbHBAXa
4LHao937/lVsy8mx6UwSJxRxOd+CSDjgnIUkSGJ/kCLt0z5L685yvm6qdaMA0IbA
VmvurhA/8aN7wRAFquXxs4+AL/rqtEPO8YahFRK7cGTdzun8aqOdWyaQxg0x/8rA
NCGI4HAxqt01eWLhkTqOtkaS7jPu1Xl7+EPG5sIEDFnmRHKzWH6bpmcyjeg9aHDv
9GN3ZO2HJ9ilfZyy6Ar/qA/cuptPzZtx9RLRFh+KJKjdS6OmdZvvFThlLGrf2Lin
cb7MEDVQguN1/dH1UToi83wQ4K2yOUDF3ZeJc/i/TKa2Ga8/cl310vfutrbKzc1g
20q5PKllknmAthcZ7sFZp1Sl+o61cl8O3rO6t01/Z5IliNT74O75P3tlbus/H5Pq
8rzOEi2aO2cCTZIUuSD605OC7yLQDJyI4J0EdCGXLC8Ed4BcV5i36MZX+vJbMg9W
Tr6Rk/G5A0F/5Nh5Ki0Q/VhHGMKRkXkMAf4cFohO6KXxS3dEa0ls6oY+z6AZjYTZ
uV/bNsr7ggxirSN3ebyamFaD3oUUqxGdy+FtN5tbF0Jl8JoH4DYQ4E7FKG9SVbxR
8phWjOfKD0lj6JQkJoDtNVScliQre5NgTqDjUsCIdjIKKqHWwEvkDPt0pW8jXhS5
YkoncIcgUkNFPTaRjHIORnPIekw4cP5XReBXpu24oRc3aYZtGdhzxu8za+b5Crhe
Ss17Rq1rtr5hMxNuZhY0rXiSWbNYryUX4A8NBQteMO4bpfqoZmh0ccZuRJZX0yi3
70bF9nQ+3wCO0upZhLw+V5bG3jH+T8rhxlBKZsICEwzj0sXAeIYJ+0YVENpnhc5r
yGuXnnG6YPMdPlrBeSwheuEU1FAfZyZe0O94fNniToGbJL2/A2ziqQWNZC4mFWxd
LPGVoWfdInQLxLVzmYJmdsHx7mBluA3kEPdF3XPJQrYtiAPfHiIPyWaZZWcgwx3o
hT2wGDP4c0UU0OyYv1GrX+5mPnBh7vfJWLdlyD2eVoVZLpcAFVqvot8IKsti8LrX
fsRiqHmnXq1lodD2oAH2AGev0kvXrvCYsezvHmDRIKocYhfZaSCZdReh2aKy+stS
Ug6fgYl54sI3tDvOOOwmVdkzf5Xi3HUlDHcQSiMmmh9oBdaKuDtp+BWDEytVkdHl
YHVKwgGYv2PUGP9Q7V40GWTbWHNihAN8zcuhj2Y/GVJvL921wTq3NMm/ckBTrRBm
V3hUeRQ39wHEniLqdsW0/o4t68DRZbtUHI3n5AvahcSQyacN2ccTa+TpU6UJqrbK
FVBDKyISWL+lWB+d4oZqVrT2b4XKqVftwqPdt4mU13DLt9/QZ8xLxAD6S6eJBopq
ECIO8TBaCk7yNm/d2Nq5Nn33Ql1G25+BrYQHXl9i1nnLPGbc+AM8t6xOLO0bS96Z
42zD3+9g10Yp1rmIgktJgYP1JXe0PCsDyEFtJC4W+HZA79Kc1Gif2p69AFDvxsTF
yURLnL6BTb34BbgzUpcBR0s48fDSqw6h0u0zp2P6O0NGf/SzoF54Eh+PfEEKREgR
V3NvsVRIgVwzFCyOCf36NUeusA469KzhTOJMymvNCGhg3o2BpWoBWI9nUohpWgkS
Yojb1GFc/OuSyY2bo8+Abw==
`pragma protect end_protected
