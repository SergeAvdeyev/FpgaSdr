// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mSBBRbvnt1Fg4xJQC1L8dKKUKw5A8trbERbdfHI1a8u3N1eNu13fC0M3rsvk7eOI
sWZp8K7GwugnHvXw93Be+2w5hrlX+/hYUyalZXjAkn0XH4FQxYv4SIyUL+qncmuq
nPcIstIPmVTlkV0F54hSGWxmVe8kozs5o25dZcthdAA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
bFiCp3H97dQm2HK6HNWwOYlEh9WAbGSGdLdPGBCK7j+WmK+vZM8RqjnufcJx6apS
U8gSNCV7N0KEKtbHAnKgIXtgq5Bi8eWWKGNlVvz5o9KFe7gr4DvNXd3oJgPDxn3i
JLUkm6SD+Z8BgqsO3CubHISgWfSzIwg9TTPJR1p4EX2b6ZW9ScI96Ztgtt02MQES
wzQjI2wCvtHl140jd7LS9JB/0odECUHI9g/+Ex5vbRS7j0zZk98YzuXXMilmx9qq
idQ4ePrjGdV+AICkMcm996188ma5N+CLN/JhUfNtvFLZtHS/RpCF+DTYkH0ZiAOI
oOIqrFieH+BQi9mbWfaPeXZKmQUje4VKC7wBUEcbWUxLVW2AxyqqoQ6eQUzYxnvE
WePjZ/oa+WCRcJ7TV2P3vhz7no3FPgudI5oB1YiWSJjAcbMJ7bJGZDItk9uprjiY
v6UDOIm90blVfIZyotaTAnd8r/FPVnpsNH0lJjnZhhNwuLUT5k3339u9iYtY8wXH
dzD5l8t0g26ord9PoidOKC4mTdMl18uWqn9FuW6vXvvKIjStalRoSd+5PUdAfFkq
NkrLSuzNfnV/ZsOcuAcQtE/OizrO0//YAkLX/TldJTtq64AZgbqLWHpr1GvV/ONP
oC+X6Qxgnu5Hjnopgq/29ujlAYL+GsOfdxb2H4nMN+q9Vsv7pYq86JrcLzvdRgD5
4klChH9Siwbyj1vvCOZHEIBIEqQThnSoiTF8lo57TrvqECqNfQ9XYk31psSxYVOH
i98lQ6iw4znRH78COp2FaHcbC3RhhdngmAeE3XXldvBLZHtd/SKhxxiW/y39p132
y5YV8r65Aest7hcN28G6cjZ/3ZAm0gLJY+X+nZXPLGbEfiW1kLA+C8nSlPht6b44
te8GUjFRnKd0azRIsnYcoi2EL4fV2wzj2Py09icrPp3PXfA6ErX5N64YptW9hBya
Pb6Epq0m/GAhByVi67xzkFP2QnUU8B4t1NGtZU1Zg6aEmzc7ci1LNrLG0kviiTC5
987s51YG8KvYLeCTTL9aZMXAHVVDKmos/OkeQq+M1e0PAjTC238QTUC5bp02RCnc
zwC6AwBx2Kf72USXQReTn6xURmUIz/LEZHK0ITV1KyDHQWOLXeE9s4pLLcCkZGAN
4usU26dPtBCVi907ObmrfK3hdaPmS9clQLvuigwCXGNJUw7QxLx011k6cNci8M/Q
Tgcdou0RAEUFD/gNxI4ay/MS2H2w3eOezGlCn9MS5FYsaTROfXIcqps4bUetdBrw
UitNLZ37ggTHOyZTAPGbPRsUGSgBcaQ6lIwNlVp8zm5Mgmx6hAM2ggeAisdFNnRs
7GwjLCQl16m4xZJKJt/4xAHvYqAOuLMNVr6imLMfmUgAl9KvXYwK2eUHLNE1RPDH
XeYI+845qf4xboM0M9fz6OFwWLZA9FaD67kDlE/l0ZBpaGFWsbKqMNexZe36wTSB
BzpHWzBAHWYwEnOpAFcVLgHwQzuVED+RvIuUmITETLpV8oWfwes+8NcrzWlviWeb
/KsCX/C1V5b+WpM07Po6zQCc9x9m1GPoOdMZNY+gXuHalz5kaetbgmvbHKanzDhV
QdcKYYwu9xqVw/sDH8cfqtFGB8g2x3MVmgAkxKOrabPDm1zZFuronhoPOExkV0zd
zgxzkc6BcTW8oIZ2jfXPSdm6EvHPeSyDrToI9l7GzuW9s44usrlR2OqAo56AXnky
XXWgAFzly8IU178rn3gJzkWqQ6rs/WbA2o1HLJ3xY2cJftwAb6Rtn7AGQkvpRjdK
+m4fXKMt5Tb/ImymGy+AfJdwfgaVlS+vr8b6OArA8ogvFcJxp1TOPwGn0JEOmDXn
sM4hrbxVk9ilz/+yFKChYEsQU/6l6u/KBg3dNLobLGoOyHYEA5e+z+Rbtb/KN5lt
v97hWKFy0AND9A4OBuA8SOzWNOihGMRky8qBgmVnxiFRCKNeb3nhnYtsO3DM7oCL
I6Zpmou0lekoMbkS+vh2L+EFDS6NVvhcqzgrXIstgKh2EiiGojcAXnFKPpd3bQOh
MGbaOyQoOC+Hqmc3bySSrn1s7XJPDpyfgpVTrtHEhGIyh7homJ5cZAPeC3EGLYJ4
2Gz+ccYjhoH0INmMPLDAJbYWc8DGgt4ONMVjeYzghZh3vL2YOWQBT3Ia8hAljeSV
BUjaIqtnPNCDk6Nw7KYGvJKl8Q3wEQLbHMp7TEpmiy5Ecmosgbfv0Utztb8dY37Q
Vec8xlYKRdOgX8m4DIJ5AvKbjiEu+j9bHp5wyt6I611vXtauo+vXF80+ojDys5F4
msSLcVZvYzCvwdTaoCah5Aj4Bd5Cb4ISxCbQXNpdLSzHm4fVyGyXTwnQuue+zKWg
QyuocG+omCtAGr89fUkuAALyojm44MGK58upfyyBoW8A8+fzZ3jj9pFwpU7RzNN8
Uex+rqk9ZBBr+yodFQmumdYe6R4qDk8+6fUhFB73yuXHIP+F7yPWe0/1KFFzoyUD
R9Q7iF9Ma1mk6GQ2az74LLy5I5clXV28LaOItlfX04ZypJtOL/lJV8fJ+xzNqy8X
GrVDBL2COhq1RWL3/GlUgPkEl2u+95NRfJgJpQJCpNaGucJKbUUKsPe+8QAyUE9O
F7dCbUhpudVgq9sLqY2Oxxgx3wxu0LenPgIYxs+B5t6MvHOvWXls5mblZqTohX/y
gU40HFS5qpveJlpoNhnANomUFrc3v0fyxcfzXC8ZpkCmFNO4I77uKSTwCaFPJJ9i
Eta9yiyr1ZEVZIKcZTQB7NLJqq+7L7zkGq47eBQ/D07MEZk26LB9cEaL6R1Zmd/x
U+9JmKvsWUDkF4ayKNEKmR661HaBLq9/U/38EwQfCzTaFSxiAJxDkpxb/MJk7uJr
EDYVpmwoEJCvQv1s3HVoCOg/Byw6sffFX6yx//gHiPq+DjwmvUGGJRQoHUsF9fhU
J70SVup0x5qehRmTVieSRwmDP9nsbBt7jANPs65SNrYS+N9l5WBtbfDLlBGj8Gut
1fDJ296ToSY0BXr53PTH8TSZGsjdr4O0/armV6Dtf9BzLMY72vqMZljN06RI4jll
yTWyAr2L/XnawOtHg/IVqm/CmUCtHRbOVe7SmPxKwhq7emE98ePD2D17hhOXWYJS
vg04+ICL+jObVBWOE70rNidfH69OnWpYWGeRhq2dyFPXup4JogG3Z0Nk7Z8Ar6+w
aKF9ukdLvN1UP81g3doCaLlqTdi+q0N1/8d/UjwFf4Nrh0bIkb6qaygmAb+rkk5X
CgPSD0NpABwhXTfsjtENuLG53Ern3HTvjIMGAnLWPTmVwGhSHB/ejx8shP5tBf02
0ILwKRMOLJV6CyYaQWg7hTOX6mUXMrzyczBsSeqeNKSvZCPtZ5rC/aBnaJpNevIa
IAcZ1pzJ2IMvmEVze+gL9j1bToymeOxrYWAxtZ5pGD5J0Pz31YOpDRyAank9/ade
UMhWGBVCDz0L7BfMq5spkYKst52qSBh/viVV8KYHocmpiR1Ary9tiupfQuxLEuR1
VwFy//hy4T+qbeOe//BTqqi4AZMlFf+z2lfZ12H3KO8/KVXdjg+xGpAnL+SAD37+
ZIE2E5z74LyFLEr0lnEkH0LjJJRyLafhaANyGP+cVekyBFD4vEvibwqNvSBih3/f
ub04wdEZTfvdQKLXlUSnyPQu66OTsqxUDG3nNoUtZSsae5REq1q+6yyzkV5JoWKt
Wk/4XYo+8yIy+8yy6ufuQvF8pzxErVFs2vCLAM84xEPczpA0mqGVoOWqy715bWdJ
Mw1kd6wHwORLlffE11DtAlS8A0QsVJk2Q/xeAP3C146hZQRZkaJCeaGGh9ghscHh
PNyVtiF37xfZ+IBeYIC12t1QfXjtMbUjioirE18bwoJL2H/KRNBoCn4zi59hGPCD
nHXV6zolOqePneJwLlPvajvwaYwLY2Es4JIMOdolmduo6kh62vqj6SDYMTi8yNqP
Zv2B6F/aAiUp0jyz6j/9OdvfRd5NsZRUX8z8Jt/G6mTEnfctN/aeASglNZdR0i1L
3XjNWeLhnTTIal4FLnPQmc3hmp9kiUBunpZDt/5VH110UiTgCN87MAWY1RsUYuZN
pmblL9GRiOG6s4hBz6rKx4IQdTBDoI+vhFJNUCK7RjgrkFLBVsx+t7zWHLTY6jiy
cDCBV2BYtd5eqypZeH4xBMawXTpDXdnY2xYqAX3O63D/FU2p9BETMz0rOlfcqj9L
4SlhL5D9NV3bm+kP81E5s38hkyMffNXWTu9Aakb/gC1+It1uHtGk56SdaX8NntVr
heO0ZGxX/hTAIe5DFOl90QXT8pe93nT/gr6iwOT9kD15J6j45zexIqZbF572SYfN
QQHQm4thf72+xYVxwKD0sblMU1njMbxgoDjYcBhHedq9KVdAQhFLboI2HNR4Plwj
2wMGyMWFLMqekw9OVG+Ve4PIdDusa2u0Zfv1/HXACBGNwHFnlOdnQooAKfG6jj6e
XaYx6yw9oY/b58qy/q/CbiiCzkFh7kXaO7TzBjN9gB5QT2LZgdXpSkTuiNLAm47e
5EGca9em+isA7BXmUKBZr/yl8Hfb1+OnotQfZPNeNdRr05HCaK6jiRhQNhRUPVvv
zOcFbk9ojzavygqmJllV1WRk1/XeZ282cNISitFc4uCHHcnINe/pnZk/n3VlC1Rk
SHkCL+5FhlfObeAQ4nUajTlkjLXQEetaGnbh3oz659hM0TIMtA9ChROwAcqWdzUC
dASljB0HCj03k2J3ss0pzmWgSKpBpzaZLiPskKFT6N01fEvo0yvkf/Ptsj4aDdm3
Nkh6t6xXshIgxUKmeqxb09wxVFsJlvsQ7zRUVU0pYEf5SGxyn8/1MsCugKc00j7E
WMfNprmofnxINqLFiikIx5c0NQqUMl99cvo7NnHOWwBXazgHPL3GvtdJq3MVo54B
x95w7d/3Ye+5tsVMG7PwUqGGom1ZnFcK8yKEEg2ZmHkU52nPQNZQMOFjphYqyIvc
ERbhVr5qtzSmnkvNHVI55wjZTqOgPZuOAUwXVycfdkG2hLWGOL4AIgAGWka2cSZo
4KnmFJD+bErWJxDKNaUljmNb/v3eN1qT0okjdQ4607cwNfUpxvsmYJu1WE2yq73K
1wioP/aqxjy3C4thGQ47WD/mH7O/hIl2/5z9X6x76BaizKfAXXFZ4c9MSG0gkyfx
2WwmXwGxVUSjj0Vhu5geK/XfwnaezE/Jl1PNVNEnbJu7JSxxxReSLk2vmf1RrEbw
Uu/P63I+z//FD/PgkZuacEmsK9mdVnrabYVaxves6jO/NQl7rU25+XBH48RMAfaX
JyX2DXTnvK2B34P8WHT4Zl2uouni+fHiz422F6O2QHvU/bE+YFECcKEgF8hWCDvz
xnrr0oynD72n3+Itrxdlw2lVBuRNWNCFl92PWEaZBfBSMsAFIufFuDmrMZH8VJv1
afdInPAk+HwQxQSTHgxnNpH7egVXEjuSfCOdyVJJoVgO885O03JC5BZxrTD3BQ0C
df+LS0DyYi7SJ7FXOe8vBmCTNfY8dHlGZtdc8h+z8neevC9l2gA2ySwwQpvhiaAZ
7sV/DcgA+NOvHy1qeUXu+P1dNngRblYV6vgH0+7nhybimUXY/45ahNTUErw1knBC
dQHAesyzFuNd0MTMuahSwW3Woczb0xdnJkqR9/FpPDatsB52rnIMZ+FLD9ecWoRD
ny02FXUfwzX6uXHzVBOrOzrPxSniR6dVGTb526nPcWNhhZB99YhZo0sW0Vx0Yj/k
q3rbTfGJG7KiT1e+Rp/gz0ayZxEEDIfGg3ia9iwBESO6CGj06B5Koe8qb+9CmUDC
b+mx5EFnLpKzLsBtsMW4qP1J1FGj2Y6uqtF45tBlIxlMqyRO96jK12iMm6xc9jG1
JbIuvnQ35HobAO6KScE9QvAkUN7F6Dw2bvcJdEsXLT+j87eJqUBasFbP8uks2XuU
M9c5AHCkybSBkS7YlB91XVig8m3D+az/sxA1PWRiD1u4DlYdqJqXXDPnJISu5fSc
nQfhvE5UyUg167rIRoDeeq960OpQKeuGXJAkOw7C+HJSEH+AJ0TWLQvt707yDG8i
gWrnBGwGFzOBksmek0tSSyC6q96apPffrQ9E6rzWTBaS9HwwYUhmKfQJZ4ObMyNJ
sCXELgWv8MAlp+X++R86oa+WBSitsI2mTJY3X3ZDEWD2+ADFFXDWYRo3rPK6UENf
NVYAgnzydxoD2CmG66lpSUSMOoC1o9Nl5hVdDLQaRPN0WzSvEIOhVr1ak4dW4RRL
HTlWz5rQgclISayl50pZK4ICffb2VgMGxt6GztbRg6OqWPsmoao1SORqXut7llo1
I6DcR+vSyhxTAD69c8Ar1W5X8AmtCAy0dhdOkUveaw+toIS+8QF8WQTTpQuKq1de
Cywf4lkEOpfoHWWSSHKMx9mvdJ0z2LA3Y2fEY06Iz5xWljOkb6/rC4JluM+nb1Rf
tRHJo6GiPQq06/Iz0BZHZbMHK5FMT8la0LhAkYWRZ93QZiPIUCwD7X7YX1pJIHVr
RzzwhejKxCWqbAlHpJqLneiFxdz7BqWlU3pbMl0/aWY8DRm9twFQ7xMPvhUaFIRf
kBrhpKqX1Gp8EsIWcp7BKgApJGKkSVfpKNaUU1llrM03qkbONbI5klmjbiOMFk9n
cL80wvWVZIcAcRs2iyQq66lM8bFFHRoyAyP1hZbZaUqxOc8M1rFrHda1epY6oG4P
M9kn540wvBioCFYrh65+U/OIMhKo6cBKjZpc/9aRXNrG0RV+g8aLMWDEvxLWeODW
TqJpPautxTrelVjumEThaSOCDqTtllAoNr7Lf6TAW1NTqq+CAfrFPkMW1fACBYBo
7LFKqr+5DY5LavcNo2NUp0G888VOF59BtViAr7GkeNxUrrLhFgdV+G8jVneXQuF/
XFHcqKsj9kOgOyKnJOK38nrpjrODPoR0WsMkaOBt19DKUWWxHeWFw4FOIuxqATQF
0RIESqqE6hSzp3d7Q/2FeZDc5PGFxh6zdS6iV1Eal5aQR9AOkn7avBGSHhLx/QFS
0r5DKKBuLx1F5CgAhzwTS3kIyDWPxN3cBm8wEBB5vjOY4kQ714bJOba6l8WePYmb
XgdtTJZP/DxWXMx7DkLyc3xt7eZs1sichYC+A/6c9TBvovL6qFybXRrWiTuIl1sX
Bb4u6YHavMuoMcSX4Rjl6AO3SevVi0ECHtloEFF39KbvhkF6/BrwYbXO0MVmv2fI
BHbEZA3ynt+1JGQ/INaHRNiVNiuH+EKIz8s+4l9SMt5aEaOumk6EO1cncgeKRwQO
ErKNcOuWpBD+HCHyllhX49TBvHLtEMio+NGmw5aQ2xaBRMfSQR/mNGryXnt7hGQt
tdcckhJwPT7q27ZeJWI3nMEgW+tssLvXRjTgW/OMChvJE8sGA/WiBPaE2RjPecBW
mhAaYbWrVov5LHLD7gd6WWnGqf7SqsyZqQ7RoeunDCoFH16h9FNiSOxS2dXnjdMX
FgiWkzol9ibMu/o1EnbTWRARBOlRzdTxFhrFoANTTWJzg5AxUCUwbcBzRUW3icdL
rG+MWI5Xm2aXGfKWVcWw/9BiHaLXlwaHYOyD45xg5bmqSXVrUYDbUyJu2DEhntaO
HW1v/RlE6HXgokeCDQoPKX82rc/xH99Hj1IL5EtsMNOmw8+ozP5sOGw2lwX13oOz
jeBUGfQjNu94IV7Z5iRZptAYXe9RZ2+RhVaFxuZwwEk68MhnHk4FHENc2oi8j6vC
0qnSl33TKauvVmMfwyNY+SkxHEd5l+bSubSTZ0HX8gQivOS1pSAk2fdwwMWoxtGz
iGVh1nzXg/2ucDMtxj2M0DvOHG1dIT3VcJ/ay//VHrtyCXp3VtE2ro3NFIUrvVwj
jmC66kKVi5K7QNhNka8J5G8OGTOOvJq88j4Lx7W44lqVCdXCbbb5ryeX0p1RgzKu
6orcfdjtNpi5DXw6v8LjQ/hsKBaO1gzTIlZkXpoEQeniBUkN9ckEVy3KCLbjwj9d
25FmOXNu9Q/MycmSBgnL1K7ZvWm5VFrn/AZuiJI0tkMQT0DhIXOBVmrkDZ2M48+q
bS3kHHnfbyVzLXysl+s3nH8Spj4sEMn3Bby0ucIcFmudjM4VeD9hNOfq4I+xPnEP
30KwCFZjM9ZqDVLQaYZ82fuj/R8/ArjXutsHi999kRpEbzwKzjjVhXzYPN93ScBO
xT08hJ98tXH0Wr0JnzFxhdrWzlp1YzhAM8JFR8NlSwSaaMBpJeCoTJwB/IifwZ1X
Lr5mI6UYHU2LDD9PU+bjSpf0xIWAT3eX8bIBFmq5yttmoyj8GKZNQ9YnrTG0uKr3
QFvPs4H/GDdaTa6AbesiQ6vSeiWmQqqxNib+0EhvbYhuAnfSb3v3Mu2Xymr3ucpC
y3HI9kb6WL30ovLfwVUZODjrlFwAf0cTvoRweh/Z0ATgtdtSL+yIFmgXUoChtlN2
Nbwpb7YyvUCFnTTZT9nc5xo8EEgiAdQ1t/cdKNy8atbXimx6dOU86f5fEmHuFa00
v8OoyVr95eJmiy7HNtDUvNzrFJPWkeB+16pwp4wFoXMPr7znglBGFjz7oVKDNbXr
RuOItsktERFW1ClPi8/vsjSeG2Xi4yxQTAzOlPKpLDWLvById+D02DR4gogxqBLA
RZe87NHIFuIHVrD7eA/KseFhLxUdqWEzw3AQmWtu3+xNIpb4ZK48yxNNM7ghn37A
hd+7aeEvj+sshHmB59bDU9YupyZxXr23Cap/k/R9S75ookPvExdA7z7piTLZJIVs
xpx1yGmsXovz8yRZJf6Xa2S6CE5eR0pSUrSWkorRcefaYKpY1SG+6k5Vqw4IELMV
Ue/bTGfvGRd96orKRRGBiiDhEcBd9Brgr3J2AWN9ji5lhVSsY56pqzMC3vAh8Hdl
WlaFFNxv7vqTtiKWHpWH2V9kNAvboIkV3zhji78T6C3k0mtVISkZ85kbMtfxXrXg
cvOSGKKEln1FDK75QOqWguRdeKib8x59knO7jxGewR5MfVAiPyJZJ8L/iGrJ7qkF
TgafxADtKfXhdQPRjv74JrG0ZdRqP57MQ6cIL2ERKdB+jOD4bUGVzvoGbhXRnS90
jHptOMTxZVXrB01pT/ccd8SN7d++ESHw7YBgr5RGL27jnJbYfRCrVGX7S3joA6Ik
vsVo9Kx8qZJ5lHByAzlNgxK1I8kpz7VFOo+ykARUcN4s3Cw3YYtvRveBH8y/bIUt
S27I4A08jiFr9Bce42ACok8VK2w9aHqC6Se2z+SMxy6+Sp4F995eRxwRMOs5hv/e
fi7qLbF06aufTRTmAHKNcTFCcMnc7xoudLGaupQ6bHdK54urcjrUjLdyLVoLKC0F
G9Ta3lI+zMRZtau7vL1F7DgOO+msTbasmAuWBYXdM+rkwM9NkRHM+gK/XT1ueXwa
Swp2nCyCDwCs5MDpWuzBAH6F6U17fEGL/L2/DgU5RjQSxJOUuUEEcteluwCieENT
bVS4khmo2PJmiP4guTbnLKnEouGblDfOmIX5+5nFtYASmgHj2foRpEQDmUoR3wtk
lYMIxBnLBuSCVJEdEahg0ZSu43AN9nKzwp/gE0XxSKik1KXu0e3JlK/kw5Qv5nSN
OmmUnig5KZlAhSb3Cg4RAS83bq0nB9J9J5HvaySazpN/QJNn/+DfrgfVsWsvXixM
QtBZUhcIYu+WbeGZef0TKBHCQxtkGbYeGWmL8ub0cNx+tQWpr/P+Cxzp719f1GDF
UY4ye3NhiYMzWd5T1ia3M6OI7Ck98MVms0mXezGiORxOeSi6ztAq4E5j/5Vk29Yb
+LzsdQAXeapeddmpMoLE7f7W87Q9qovFJyTBvvXqtM6gIesk0+62k6V9huqepqyf
X2VKLvhgRKSM+3dQSjOX+qT9WNDZoZrpcwavhPHca0wgzMUB8o/rjvPqYrhrJS6E
sKPrWJLSB2pnwjWdQwOSMafpj35nx9xhUNSnAseADbgeeOdQ9XiWlxa/zcriSsGY
refgCILggM0wxSbktzsqMnuBlM+tqqFIB4SJy+CoyLXYGbHO/AWKAJFfzWtk9OhR
vbgr8ZhwfE2cnzILif44p6RpEQC0kfLrRx7qiGY93Q7PdluTiR/77DwmRl4VITAR
3EFXD0FL5dh7Sj1LHXLWdvEZcwP2O1dfgfgcDCWkAgM6NFG0/ONV053DGvSbGlnB
txaObKhFeCHgTNZxkohAjkcvCXTb8jH6axauKesGEAjrYVfIEB8IxpZFstCgrqbB
5qWXDj0l6uNW1o8fKpjPyMw/k7VBTl/yPU7IGsmYntoFOc+WIlTbvI598iFjU0rZ
vVQjXX20vkYFPwmL20YbD7I0OlR8xAuvkhe6AZqlSgqV2Yuk91dFfKUTz0twidh+
jOvmUou0Uli8QBMj+Egcz+a/zYpzlSuFgXBOf+J7tyiYrG+OZpgnnSBSaMk0R3Y9
PMNXoF4Bh0F5lZYssxCykyr8Lzr34QyyD1L/qLDYfavDnVmhIF0yqY08DHK0Vwu1
V64BzhyUimpE2RWJ0YFbfS2gEuvr+4WIKSBLA973AwC+lENI+mviaoMOde2leM+r
XmBtGeeqFWOhYqm7maXiyq7WANf3S56KhiwZJeLI02VPbPq24BYmORpfbBENSZkV
cu48zUNdh3ekkiEQDO1xH8ER81AwVic7/LM7JPoR7rue9RN4+C4YwSyFWK0TD2Bb
kWsu/BAf7ES/fuxNTdrvVl3vEfDT2rz/TlGPN20d50gWYIz+B8nnxarXo1OI47Cu
r3jVx3ZmubQnevjWZFfi7dg0zsuSQOYS9851wW1ovLn9VsyQPxGvm1dmZCHgwrRd
iBj4HckhXS8mi8iFTyPALaj7SNfhTEhiA7b9AU2xKovBpCkRKqoGW10DU3GLGJMj
Y8BGrzcz45iWDiqD7MNdskEwZEs0uEjDlKi6+NHFX74u7sGozWH1jWS3qXQ9Ia4e
3BUFYhC02wXjQU/GiyQSYN4Jmsl2l7Bq/7rrObpyJVzhRKfeSrxn+I10NXMbehIx
csJY4zZhTIO9WZ/vrwHP5CwtOBDfLolKxVTQit6lUK3nE3m0iijYVpBSUnyNi99O
A4zwV7R++4bfaoaHCBBzrRvWRi59NK2Jp8h6fOF/yTUKm9bIyhyOvKc0zCYV6FOJ
H5hW7q5dfFcZkGqp68P7CZHfcQJmgwA3kJfymzmA+V/mT/z40GvkFsJfbjGbRD4Z
hEYIhicXu4sW1hmx7VKiWMG51OnH6ZUb8qOZckCPfovyS1QvHkoc12kfVSz00cU4
YzzVpdF1qs3MVWVSGxzW+1QFJ5TkS561raM8xoOJMrERv7OPNbnFj0wui5QxoC7z
2gz3VDNgAUkqfdOzsFOfECVIrwcfKpu7BAdfHQKASab1a69UnrjXxHt83RZ2Mfjp
BCigwl+uuhKIxVjOC9lL9diJ9Oa+7yfEKVX3YaWKdPTttf0JE8OFXm7xiAZIzYxk
hTpNKNdaa+S9pD+i/dDHYtap8cCQpfub0TIvHEUJ5R2P/W/VFwhU3EgqQ8FCKINe
bnD4mQZk926PMP3IVGgafzyvxp/BZrMQvH+iv9K0D6K+jTQcZ53/8LHMAsOsQfyr
VdfteT6p0OP4GtwUDj3Zy3fzLAndKqfovnV9rKXTJTjl7UydOO/QCcY9NsQIdT1+
1q1kG5N3GjG7FB/anMhnYMsuXOx440paUdl+lgKDt5Vw5W4RpfJ0qozXyBIu0aB/
1w6dxVuzvIvtSqF4nE3QRXgbmInUcf/8bNhJ2GEa1QwtZE7UpPQAMrs47XonSae6
tDxnF6NJkVbWQNdbIYwA55Yg2y5D4+1f61x28LMvTaEhcl83Gv7fOITcmHAM43vE
DdYxeIaQ4FAZAzC9HaASVUZYnXkb5bFL6HfvvXDQC6LAO5MZA3NZSlIBZoBLdQWU
9cZvUC9pnro2emRIHqus1noyAQSYDppzFLJ9KH5xnS+AgLpVeaPZyvUgywU+9R5R
7isT2QYR/NSB9oGdzcq8yQ5u40x3dgprttiFvAiKuzFf51IWWwceRyzHQjnVSC3e
mwEaKcPhzO0Glbm1JE2nrq5e98c6JKoIRe6iO8aG3Zc3k/9DcHMTZWRBHhdJYeon
nvKqTfRnfsREioNa8XANlf305MKMM0jLb6XCBOkP3xrT9ob5hfzs/so0IwbQtdc1
hfF/IcxKiPhFAEtn2cjnUFQ57OcwyDGhx1bgzcPLnafEunHFbcZGnWkdnbCfYzbJ
vQ6//zKi8u3aAFR49cLEO1Yg7DDWPUDGuR8cQu8Xi74xARk9DOSVbyDA/Zoy6dKh
tO4Lt5r1uMCr2rXdWlbihzCeDDsb77ZeEgi5sDQ3EREYqQCVe8j9twwFyji+LA2j
3/UpreSfFSicJ6FLuGokf42akT6icRzx+FCMuLCVTmDXVI31ef38ypLUiG4M5UOH
WiFxv/SQSQF2bmaTviP+2g/JoSmYnEdi+ZYhN73mhOsPbHIapLLPZU6INzts9zHU
RUWVnP86/WjiPmPHZfXsAuOfALX6wNoz8/5krB5KS4sgC2OkmrxToCdxjpZPMLg4
gwAKY/zNw06pclVkVG34eEbqkYfkuFBm1ykFoD3wm+n8b40H8OmtYltqbrBiuNx7
c1jP+9+L1C03NNUgRhMRXeJuOsYA03U73FwR5JAIBQSe1LzR0iiBavNaeheLDKeb
65jAQZPUiv94TGLormdS3pxMKiLZX5w7KCJ9PWiOCF/NZuaUIZ30atdHUw3VP8Wq
d8IebSg1RF+TT0s1Bb87lvzKpYnVonU8Yxsjpc8Md3rc0MFH6PiwTPBMzVufXhyd
WJTP3oMa6hI69yPUDg3NGZ5gQXSKX9jDCLVNceMXUHBF//sB3QAZIYKJgUuZTAJ2
ZLrrYUv5bGLIM3BjMahvPjJwMTc0iOexDcfcFMx3SYe9xzcAi6WJBpICLoMYw5N7
nE82EesZVkhB4CW750zORB1kKgvuheAHjD02jE7Hg4O5Eu6ukcbpgSn4v7YRRNDp
RI+j7prVZGcUtJDpP2JSD9koL9bHDhdUxV+xiclRApl2EffGNOMnWDhzP5Y2yxQt
+vOfyYS+Ujx8NRK2MjiSjv+FJgqwU1Fe4AXbG8cjEo00miBUyAwBqBIr8+IY/eHU
tfTaO1T0WjQeVdgkvkuMXR/ZXtVvJN2vv2JZq9faiH6//YDm4RuPcwuXtOh+8WhF
2XWJWld6SIrl/JGDA5DqFacbWk+UtaAaiT8YsfR11PMyNhSoJy4Yjip1e5/eU9gT
Q8NfQJEQ1gIKKHNjt/3Gv/f8lBPqm+vGHM9F+T5z+qKxeI8EhBltkVUF+nX0BLHE
NKZXrr18tG4MavNDgtlfi/oK9O5HkOXKr/NA1c57Q9fNLZsOm2OSVY3l92rJCg98
hClVzv5QnYEnjsobo7mMYIod+ESZd4WzK4JPWfa9t6fWMPdT+GtN9i5AWfK1mVcm
v58Oq1G1+CCIb3VEkgkGis30pys31KEFPlY2illaiMBBA4YRfIlcK9GDL19vQKke
nBsV9Fj9OKY5QXIoXDS/vsP4rhVfAwLaKyyObT3DAzDGhY5wNVhNU1w80rs55Sf/
8zF5LsJUFWxn5ZfNlozlJ07+cVuL4n0pK72umlOMMoA4SAUe7SsS2wRw9VEOCTbi
g3K7Ck28kiZmdEQhQJ9fAlnD2C9OKp7yqXN1lZMdQ5WN7kAbs8EqUGhU5nw96bb/
fHHBJo/lGFf1N06LcdHUBarQgw7fQTGDyLbisMHl5HXsS6TRolBSw1KNtYIgmbGn
0oWipbXUqtSsUXIG+HEPbVsEWrT5MxoZM+1JXBi/ytUNLMKtQTYgE+q/EO7f2ad8
rkyasuMqpiMLEVuBR5YJDmkK3Ii01cdjPELfRFtGW1GcjDM5W70W2DhvVbFZ+rQD
DtAR3kO21TLrvWSnGk7DETyASWPsUhMUQrXRPZm01vxzpaY6Ou5ymFD3fX65GHLE
W6z8IMv/C7zgGqc2lTJGgC38f4VkYuHaOGhd0qHGLQU6rgoBYCLLwbLlMT0KNvY/
+yAngBmZuXJarS3rKG5SmDNbTw9LQ3D1vqw1YkUHS6rGEPSZIvemfkdkMaWx9/sB
FYZbgjHlygNGKDKZQfHOpEbAG3TZAniufVe5ujrqLoE73yzgWZVNiH225VUsuWnY
6Jif8h96MaOWoUADb42af4hPos+8j8zVZKDoGtAN6q60siLt3+Uvxbp9rUfNR/Nb
q8XvOhEQCRkvF7hoGUPxC4Idt1h0HyN8aii0y5dHakeCgsEyXbXfIMREao10Sjyd
WGe3uL+nzsuuCDI1xT5HazB0d5dAI0kL/IGHjcZQJ7hCmZWlLLJXgZI3lvpOWPx9
h7Nrdr96VTKVJ2SeojYd2VyKOj1/4A88SSYJvtXzUOck/675smVUX+xdweQtx5aw
uWO9Wgu4fYb7V2+XqCmxsmt0BbksxcRo5Ya9nOHPWom+y+ViJrqbdztjKLufpko2
eDfL7BDJRoR18yWyvpyDRI7IOs9JNyEDzE7ogN50PDx71FvN7me1pS+nW0LzOlOk
eH3/8OGBEG44C68uoGCrRZFf+MNoBhtJpJelprXU0GA8CkpX3YffUV4E6ftUDiTW
ewEwtw6lCrsrCS8pvb1h7nK6Fb+AQ+9W9zUIT3a166Tlud4Ez1/RN8bg2pmZSn+g
/6VHbeJclEGo57Kx6rrASJXY1OxcsWDPQbEurz0kVQW+oTaZtYZJclRB6fyiUXt/
jR4nkb+r80Q/LKUApLvwrLY8z/Ygk04MRT2n7bAzlINaEQ7etWOjTxVjlNvTT72v
qi8FB2rITD0/90GXBb6+p8CQvot07/Id9eg1499roMcqasp5XXZvj0wuSx2DbA3y
nXXrZXxy8Z8Sl46kvpz9iB0piRV5c0fW6LkqqKzhRd/gKn1WCs2e+7PzEC2zPFjp
Ktkgx7kRlVr3Pn9znO6NdRT1U1WRYyJzM/W/KsjdAHMCrikrPoBWN7kMrLkAe3Rn
QOWWIU9C4/g4Qfye/zACnMNQUIInys5usMJ83YW37fwabcOhB/vBbZ/ps33+cfdY
HebW6iaZhdv+yJISXJVua/4SQeGiY4M970TSs1ifTEkBQxfbi8S+20pCG0SFqAot
0nYwEt6Rtu4iyLWQPVdzKNob2j8yWfB1SQmSvxjCpQg2MAnGJ1q7XgjYG8JvXIri
zqiMSb+r0W9HGm89iV3h969418IGm0SZp6nMn79kvl7hIy2xzaHqIXOICzGBlNuT
bTm2pWoV7gz/KQafK2iIh1TRx9duytdGcjXW9ZEJ1e/gO37qoFn8dlyF2QUoPcAk
W9SEkL8I/Qnp2I58O4yFx+f2R6wayQshNhqEmAwAoS1WSXCs9asoV3PZubrIyZ+6
mVFVcmXlhKChGDfAfI4BWV2LV6K+lNcA+kKcrfWI4wZci8ysTImI8xZvKhiH/GyG
LiGzR0RXK1oeoK2unU9fagvYsjjzmOhKLGyiqsoKxf83lie6+2vAno+j5d4diDNR
9uwbDr91MRtxT5EN1egafciH1tvN46Alah3L8MmlM7FZZcr1iKGGc46ayTb/Bu1c
F/V6mNqKyXoizdLJqDXWHb9/PDEe/4YGB8F1yy2iMTM+VnNML+JFAQX0mkm4f2n3
wl+Nx/1JLnRg20RY1V3qI2hQRWFpZiBEar6YkygYqyksiDTIismPy6I9zYS5VWqO
qAA29BzHAgiUQ3LYZv0h2Rp6MK4GhodUNTnLVeuv52VG9l4FKHETyKAEzEH99eUf
QPWxk/3GnpgQL13EIEFu/Bm9Y87hO+1tDqEAyzctcDbIEd3fE99etuSGlxPBMb6C
Zn35tYP1x30sbe/QCq+2hZbNiWrhgTJ1sP7AxcnKXxnXL5XEp3oQ42ILJ1ToQzP5
FZif4/lUp8trr0AYiImYxt+cMhBQfm8BJJFHi+S6wrIKwYSsEDHOU/mwZ/i3ee3U
XNb4OZUp1b+LkQoo2yjbYKfkL+tdTICuS2/3Lux2KFn2Rvjq02kAt7xh8zirT+jl
wPU9ewD0qOvuHQf6fiTx5FduV7IBf4R0C99gwkO+OdTTHkboX22ECXxb2D8i1CCL
ScHakFUJv39Sdxga7LffuvnWaWtZ2kaMLYVhenNk1xbpD3Y/RFyWSSmcKe0OEu1k
O8dm3xbYgVroToCQYGLct1kXrXRhp+/KetMhEbwYctAdBMC0ci42NHiYqlMuI4lS
2LJlIqRn4IDEIpdm6CbubWQU98RpoWnh0D+wmINcB/XJEa+jTYFP6RbrgmNS+atL
sNsV4ITPLs1enpC2KNCGqCdxpBblEsDjcuZzFVzZZDuh9JYM/LAG6csM6uVB/Ul6
uokIWeSxR/dJQ67EIL4YKX3y9ceKMoTxsdAJKFtMmTZmIUljNrraQl/PSSlTK9Pu
FUUXTSSQbFsf0r/wclBukVSvaC4XBf2XJLMdjN8YLRjiY1uWHTf3BADQx/wjdTIo
0SKlHcxeWug8g7we8hWJKAgWCuS2GMjVj3aP5aG3xTs5CNVUYS5N/7MDdNs2GYmt
nrv6DECK2ioSVqiu4PkOkgFVCRHT/Eqc0G7n/fgmGV7ltzMNeF7jAT8VtgkZ6Ed/
B5jIEDMPRZXow88VlJtrPSnNj7YGVyc3f1HvIlkyQIn/y2gnzYkWkvrrrqmNEFqS
k3cHmuUWaaFTxSZcgCL2ipPknjxq+t1pH5lVlV0y3PUu1MOGsoPTaZ47rmgfXZQq
ak8IRmw2eWxPQOLXbEkVzfnZozF3mq+zsKXTN/Wau8ymY0Qndw+4VLP/2PlQoB6c
l4F3DUcuHVFCKauKsRGDgAPvxa6anRHbyi8pCLM3HsEGyfbLXmmJIxWEG6fbl85a
Q5d34GiNV/hjfnXwDmpBuqj2dVaQCYjB0fw797TSEumPyacetn2VP2VxxqCgI4tI
+gNHDodjtP1BaH3KD7IucNuuUc3ibsGnqV0aQWbSrwFAE+57UTeqbTe0nVaBQaih
xhOTYQZaFJo62RS/7PRcnhOdnz44c3gmCeSeGeWTomBJtkUIc5daW16GcInOjstJ
n+17xnCCEBUeGbC+kNbKiTC4TFBXbSEQ7uUpRoMROXIS++AcPmIjxWhYtdGJxs9H
4eodp+cDbDFT4SOhQSS30TwQ/ixM/8VYDW/9g/2wh/S5mjhuh/UxMZ8zGBn8eXv0
kg8iUqieAz/dMEr4shIgwaRaLCpzQvr2zHmNuprQPhUa8IALtC8Cvvg/rWqfpsBe
5xzKoDZOJcTs2DFzY5a5MYJwuvzzEZCCFFU/ap7pOoqlUhQA0Al+rHAcHwThK2+x
+crGrDl7ajPT69UiAfDp197Zu2JIcbe62YdjsZdQd3c3WrEztlrmtwv660Y5dKmG
niV3qS5ZM3AVvktS2tZrzgAINdPh5I9X/xp5+hDFbsJC3M69FnAAXLUQwyn9XaA2
6XVTmMlw/3ISqr8ZWh4Wa5Kr2t6X52/z3loKiwsLzgTgw6Drf0rlljVRaQjQb4zD
uXHrZzZjMIflGI9Mf1C+rih0d2KXgnXlKvwOm9AL9ZbrgBPcwC2ljEjbf0YyzcXF
mSFewLohGkg9diVlVGwGDDRC8GQ8qVDONJafaz29VG1PHVJ5ImAs5qzkgfMxogsi
dgZ328sSjwnloFOjZF58cY4g3H65S0XvFsElTQB4o0gkUN7vgNnalmDzkf2CWbcJ
NZAq/bnPmQgZk8mnJMg2ffCacTM2vSQ49wuQ3iKg95PZt3gP1JARpN5CQX+aHH/6
cBqkJXplZbPgBdnhOCaMn97X1+O3CzmrNx0T0FuMwTQ2QjmIq3tUdxD9Tit+dMt9
BmjIbdEb2Qxe367YOw1UVY9fFhA3P8OYPOOeex1x7eLB3C29SpF6Hh6SpbiibCwC
cnEK46ojuGuGurEBhS00cj7d8EPh+tHUg17/jZC8Muzd2VjIs+7GjTHlBjyrNML/
EpcjroE1Q01aepTPbreDAGvRf1XvILj3r+VoWo0tM9TtlBUeE436c3Yhk3jycs5J
XOrIDbzLB45LBbX2tO5H5oKYKQqTw1NZIZ0Xo9ak0g90hlvakYcUCM1q45fBugTw
2GX1LQjzE4GDhM6BrlZe5uaaF8BGpIWnxdbkwUrnh+4JUUnQ7lsCti4oJXzi2YgT
A58dQcCJeJBGzY6yNcr7OzTf560h7kSiwQsQLbGMWA41ymC2MX28KIl99zfUnL8C
I2n9H6UGRBDJkTqKc1vqOGfVPwB7bImS2XBLiiqtWYGehvMPYYhdTIYC95Z7Mre0
D7zCuwjnoWgk2BlDDD3dQlzm+NsZBt7p4OP/sJuZpTdfg6idngkkHEMgHUZlNyn7
wBrDt0mcdNSYfEV8Ge2ZZguAMM/rj4Ug7NKAPhRTVXntJduENyABZj8g64lgzGSo
NPMwQyLfSpHmKCVqKt5wLqozzYTcJHEPrmZJjMcAGmvcwXoIVh5NFGbQnx8ULP5O
1lU7TMOVunKjsim+oI7tAPNjTE81sbLeOriqjRIcKqDxwZCVH4jqTn6lG17wHYkl
seD3Ha4ZZ4naRSiL6z4J3r1U+ipFjy8sJOXiZUSAOtyaAitxxIT2K/rt/o28O8ch
dYvwxkJD8YvIltOLhuUrpP1QjL6hVHy7UOnJxEJlRuLjyg2RO7RzHP1kib8dQ2vE
3Ki7Eh09a+jh8CN/H+xqJPKhCwthE/vE6NxBEVcAceEva2vUN+cORyOROKg1hwoI
qZ4JBcFnCHlzG+DpOBchzxHJ7MN/Fxl5IgfuUC9DaumSPP+RTvXCeD2N7NQZdrN1
forIWYc31KQc3cu/ZHQacw==
`pragma protect end_protected
