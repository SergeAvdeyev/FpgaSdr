// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
t/KYHIxBJKHp/3on8/AWjhnM0WtXtFmiwrO1qr2+EYTXgX97vK0d0Xr+7c3DEDTaP7ESbBKm7qot
YRpF2+4kTzm71BTIkJA1AmK1M3forZUKZmkbL7tEf5QgANnDoP9KQTlPBHd67N97N04lYfHoXvqS
GIsJn9M90XyGTib6vWGr5YcPApAE9qp0fyVPjwxBKAKk5UEh1dtEaFQWBJQr6pW3wNzXd8VJ9aZt
EafzNSVEeeaVtrctBc3AwXF41Gvm408zDyYz9JBHWQdeD6v2qbYoMm2K1laPcvjKSRctVRFrpKRQ
mlUPWLfxRwiOZ+wTkAeY+EQwLiLk6RrZN5BojA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
nxACube4o5uKrvb/8tM5OcMU0SkUXWg/15ow6CPT8xiVysyxcf6E5uBhBUzrQ5v26bWm/M089QF+
Y7oU7NdONHBVFMGEahR914HD+Pc8pm8bQn6uDLwl7fZeV1Yg98MYLsurNcbpHcXE2Vsl6kZXR/5S
IXYbSQvRHafeP8yj90SFDcDOWHECbZlsLO5zumLRE2KKBkTT1iIQfw/jDPOdVnyiY0aKrGttdBKj
+xIL0/HxNekr1uJ7B7LSg9SsMLLgWNU/nwa8t4KoVGcuAeuB/q8mgbinrjKvxitMYoTUADrnuOvu
u6u1frpvys1f4bOUKqa939MEqpRFJShFMfCc1Js72fUX0yxNA89dI27P9E5D3hFH5QMLEueCJcbT
s8uHHJWifQE3YxRav7B7kK7laHVuHn2fsjhuiE/PbrsYDg5xNMNmZdhzvDTk7CM832E6VpRB++0j
ktI5RQwVTqewPaF140NaLOQ7OPaRqQ7EGC9qLROlIToM08F0GhgQAwEe6aGxLecvzxJ2h6A5/FtE
u2fhzwOcpw8wCW43gBP+mLMI7bC1MErw2SfTZPbpAdWBJFRcJotQDxPtv5JnkMgOCZVVkTUvfY62
0QdHWazahwhTFnxDHPk0UI886UDFxQ74nqktPtM51+uUV83VH8D6jvOhCDceC+av+e/3RDYvVrPk
BUFfeacNGmk/uTyy17OvQEBiH37KM2GwMS42+h8E7gXbNuIpr94MlF+4x0NP7JrIg7tymKwNpSEB
SyjZXal8U4hSaAkDh25kpofymq8Dj+JzXnL1pXB5jC0VMRSltvQAVuigZiXv3w9OqCpnmQZnvNy+
Wb2aRK9a3bqNuGL8JxSC/HURP6tbPdSTclMIUqLyQRJGWLnWDoyY/69d2eCYumBB2Vm1EZcY3dpK
g44MeTv6bN3qfGaPxay2n6+cX37W+7tASS4j4YjPOLhpXYy55f7WNPpJqbW/+vPi2V51V5x/pkDE
kLIFKsj6yQ34a3fLuMcrbgeF46LPlBCrAkfgbrGxafWMGvWpb3jdwNPMGtJmeRnSgvPd3Zm7Wlmp
B//KroVQbDXqWli0PAJsJRoIz5Izma6H1mJ3PzSCV8feAYiROBHiba23r9y7RLFTnF0y5H4a0fgA
YEmSnWlcvMz3MLIbxTCdXOF92e50ExXigZx2d2JKyo/SlLU/Fgkr0l42rcWeF9mma77TRrHsZajv
Hcd6OT7fMo9XdenDWrXmoo++zqxIHJKf5vMBQOeVvY2xHxRUTHMW5ONPsyVBrj6LkLFX2sa3DO3m
VocHSz5XpqLq68c/KgaQbfqPFFMT0Uw3FxJTyCUAYrhosi+7rimGjAFuOrRaeZSiDe13AS3v9/GZ
4efjwb1FOOxQoVGqm9WQ1dRRDIbJ63fjnJNs5uSzeHPFUN/uiOgLrOi89NvHT3tspNAw9xALDnWb
Oj0cdgArVM4HK5wdVZIBDqrBGJx7dzWq+nOpY/nk0Iy8iP5spaMY5Z8F+dD2muLOopOxrDmmT6KV
rBxzyjYDIjW71+Mcmi9jyggQxnV/7KqYp4OCeqxIhi+WGDYBjezCfJSTo62MQztPUO68b3PpBgAe
2t9LEijkqi20k+hHBL9HTulScy1EMhX3cUzWi1sApRkoXMj1o7I7kMaLK22zQZ2Ku+KF8VTToJEN
VCxHLAX516g4cdtR5QK40ESFHv88+fzYG6Vm7kOui5Qwzb1yzQnukj6Ez27u+BdrO53iWBt1Zw5t
jxndNZlXAOMs4TKZ/azxgS3EsGCxpsf5BkI4jP0tnVe9IGHSFVTwwcZH20nxYUlk58nl3M8mDs1Z
OKXsC5lrPbJ3lUlJybqo3hyuVwZpRz5GqyIjXrmstRBRxswELuv9Cv275RHsqJDsw7H7STWCX2oI
lE26xNW/r1avb0AAjOH3Ns3nmyfPtyUhusXf/ElJyygGs5ECo6uL515pwdwNE7cgNsubA0x3X9KR
A5/9ZLC1LiEKwYwp8JAAB2XtEoD8FFI0nC2o4qk9iyBpRfm2w/azzFaW/eoEaNtifhlAj27jluWQ
iViYJuFjJ9mksRHzyzOPQwziSkw3W3Wdc76O2LRJk+c4d1Gf7jR2bC6jmmQGj+8UKZR3hhyqyL9F
2dB+p2mv80UL4tJo9qZK4RxvVyMxzndUFc3bSIvqH2a4MWsem1CR8FBrurSJvXteb5vo6ZlX1yJr
x8FieprP9yKMvwpqCerWJtUom/uKk3gBc2ISf9aujfNvTiVbVr7h+DO9MnKASWoeoJlEXATe6ZwW
NWZDUbDY9NxnUuyslwa27XIeLhavw/2Qo748DS55AD5PHSkcgI5usTYqouyqGyVrm93XYfq3zEUt
PGtYQ9ouBgtu3zUPR4LDwJ13hmB2OC7DrgkLOiXXM3cBriwjDJZX0uD09ZuiPojXA2ZgzJMMhcer
D0pNYebEdnnVTI+vcIaoUqXeL9Gfmw0tBRDqhti1xbDZj7A97gMoM9i4wnax4EGjvAFPz/Pugj5+
TgrU+HSGLBDEDcVRsVP5w6qSZSG4k4sO0JQtZvcbwT+Au+gbuNhSsE1tLMhx7Hg6Pp5X7IN9hcm7
yqF7lVM1CxYz+G1NOyuN//1/VWAC2RUsLhCua2x1fz8Mh0QbpLc0LJnaTFhy13McamWl/e5BZHMG
rtmeCA62ZufOZQFo5xMlIFUiUnbOP3I6elFzQeh9iY5GsLML2SoGJBoRG9NE9EF1mOE4L/MCiLA3
6Ia9+97Ikah/2chLrT/GgGnpoH/hAWIqaHPpRp9JNoQfwqHg1DfkDKRsL6ekFMoY0Y1fPmOgWga4
Wnoa6TZYHuxV5E/93fU3Ivw7pXIL2R1gv6NQWKXviODzUduu2eX8FOxEvQrmGAfkHvnr/h637mM8
NcWjJSv8rOEs8M2A+dNmhRoOlWq/kAhzfeAb49C+oJ0xBAEo4kDbsp1l/dk/UXxvKCaNjpay/wYE
dWint5K5jSG951ZdT2wN+TZJRzSdMxlx/RGtvI8CvrA5gxDSW0ewqqliK1pyEwVBqM4y4WXZ7vsK
LGj9+y5OIejjICm9YqKrZWSPyN5pDSyjaoGC0+dMke9SvofmF+70vvrWqnOX3XHhx2B8n0owUTZs
QMkQLCPrOvE/BTQ/QtpHHG99eqTv4IY2CccSiPhBdjx0KZnRjhYLxW5kYo2Z9s9zGYwBbzTGqYlA
Q3hDNSy4YBI7UWNfzlKOMykGCm9Rn/jkBxji5HXsaqQJPZ8Z3MuszSTHK0m8JoAd8qlEfzhdZ5ub
0jtnr6JA0GGXVKTJkB2Prr43k1EQqLiUvYdWJa0b/A7A/HIkBqZyTzU57H2tgK687V5iQH3l14x/
YEvqkDLcOgfo5xIr2opQsbRdVNkYnX7hfGqbrOTB2lNT2UZ1GS5UcPBqikQEY8ZmIG7rAJR2LNev
2G8635UtpnpGEFDGRJRqYH5DGlyJX01LmfPAtxUd58DC7tG5iui8HlYm+8v1jykZSqFaEKN+UoHI
workGUi142idKDK/VO085axtVyAQILPBk/tR7C6w3tHyf3413sOSs9FSXvqImEbH3uhuNGuDW14u
2Gw9DMt2lRd9tRPplWjqynuV8XgR0DyMfGsC1on5JYNGen0lXLV+vIzytESeZsg59HES8GcZInpI
mrg8zhpJJ+anlTgjxte30yfUOpYjSAECc13/h2QtX/GHHeapbU7ENnA7LWgPgjYoav9Lp1ALGYNy
GDM7D4p1yn4IIddbRXXFH4wyS6LcvKA2doBrqYAkvEx/ZvTqhH+Bjmb/ylgqCY7LC9cclU7+6q22
LUvNXzjr8a+k8J8xiqN+mKHRl/JE3C/jmeFtm6yc5QIm6U1zXJ17bgTys6C3sO8ZnjRBLNPjdu44
4N4vl5o7kcsnFkff/VDltijk3UiXiv7fAnStVFT0CWlW7zijouOA/48XlF6Zb45r8Gssr2FkSck5
wMya0ke6cauyPCmFQjxvSf5mjVUh6aszbWXdtci3oBdpi9BezcAShVGSN0p87svSGOATZqgBrKaF
ogeiDEftA3QO4RK0hI2pFfUq8s+G2Cyl34KtKFEGjTxqu+cvyYtpDt0cTJMpEOfqTxhqDDrh2nex
MHn0a8eMdfgRTdv3nL1n3B85JYeJxUoFuID9pAXwWMAxH+STUmJkZ/Jaa1X+5+eBmqaD9W5VNpI5
+KmPm8Bf2A6w8dYgJ5ssclAmmgHpfWay6vvrZ6RigQMFjNzr6jY5EBMWIvuUwQjerqzUcYLevmpy
rfDGykswD9GVqiteCfrrJw6cZEr442mvvHOl5WxHh0T+OOk3FuOm35JuSWJCf2PUW9VTL9vlF2b8
CU5aAKwQnJ3NN5/xE8laIPK1b3Ogv3p+Q9dTQ/sP7iYOBtPVfCLSbvTNUeQg5OH8++KMnyF6bee7
JPEreJVrnYv2X6guuKEVSRkQEH6cK08C+Fkefekv86aEl/8CHwmy7W4GhgGxI2TVsl7yGACbtrSk
df/MuZokiIFxi0b6iDCWgnCZECiuH+5RSCSIBGeEL1s0ibfDJopWJtpkmH1ZYCQzuZP1IRVxhbIl
LDyUr1lU59mvnipLiKMSr0+HeXrKv4znEU/R0nOCkSzTUiZDy1k4o0ge5u984C+4FXIdk3F263lV
KytclXeVBCJgb9DPu5wz3lNFQ4wHdeuUnHZve+LnFzhiuYcmSPW9bmo+Duhj9+Iqs3yfcZB5R0Ue
ps2Pxk+4TEuYvPPVBOtIDNyUB1djk2evYbBymSDSkt39doEmvCUcGcAtVMqr5FH78KQXtvb+Gxsk
XLUiMq5e7tyO+7l5rdZeoipGTIyKVs88+USf1JvGmMQdnSLn7qDzAtDQm0lxBK+VIDg+TfqIRE6k
6ymeoNBIpBbW6NeiK5qHBzXjAZ1y+5WI2/dobduXrRknyFQl9MWUqFDbvaMMDTCnQb7YB1SlXOPa
ua7d1oKhAQW9+g3Al3lAUneb+PMDNyrxyKvF/P/5n+HCqTxBK+2FkrWvFsa1FgzY/E81GaD7tLIc
/cuz465zW5v/T1OgKjVYBKOpuJO4DkFJ4QEE42D7Z2bTg9I/NQ6euQpTtLG5+uxkcq/l+3JgNZdP
3elKH9hsSFZWJWY5ODBxegwOwgto0ogFc6VsbKsGwX63Pg+V2GbQBCXZkrN4lyjtGAZtm2hxmnTW
evjNB1Nv6+Q8v5KH6vwuh2j01lOnhY7wNz4DuAi8TXtCKw7LbQklK1tS7WOZf9ijo0u4ehBdjNTe
IVxlnadufIWRGb5syG8ooJM8miUIQg+Y5H3wubg+HVaErluuJ2LkmnDiCqa/62uPI1/IVM71bcWA
NhGvzxEUYYb0UNmV/ucwyOPLpxsriUve4xtrwZewh52fL2FDedci/v5N2YgVz9gJuh5AZsSVJO8H
KK+oeZoXoRK2uwGfF5aIQtkSO3w49z0oqocrFyyRIENvJqlUMxMYLJVkHCWT2mPPpW/+4BDlda4z
mkkTE0fr2MUpmb0pdgcQziQQxCuENcSbUln76aEUriXXjUhy7Qb0SY2+1nFOygjAovYS3fe+D2ca
Wz03Cy1ubx2CGNQG3JKwqtnhuTo4JpcYzcmur30XZYVW+bzgw7fJwcsIqEUGhjioKlOpJTrxMagw
9eLceCvWujeH3Dt40Z/PNwF6rKaYnP5SpjcFEiH8J5t+wNzTJwajTEyXm/AD1Hksu7RjpbsPIehr
JkCzFzjo6F4IBSCAnEqwoNg7P5MzDDio43Bn8CYWZ0k/oYJw2ftqe1aH72X58GRGE6UkD6g82bco
fTfgkjiAWR2TsOgs81bHgGIGr1Zgydu/l/p1Y1Lu3Lld1NLwThSnm2h2nXXhD+pUs5XNv33D67Wz
TFb2Rm1lj09gxgtL/ce5Ww0j9/cR0EOGrJ6D6TCTmXZLh8PfKmlsae91vQlqDylUfSOHLex1tbUz
i0t5OMmRql5b9JH/Y9CKvj7tZjjVLhnOr7Awoq3lvlFEdhgCPiBBu54ClvM4PhaGKzwuk6kv6HzX
n7ex2zamntgavJSRbebnS28+ceCWE96I/v558FYhjSwp7cMWr4DspNJcMHooGwWUNoGMNHg/3thz
cUPJRiw4g7K0m8oML6/ZC6Ae8adINJgZ42386er1CRuERRzNTqm5BJvrhIp/Ho2BqcaWzOMvBaY7
Zv5KwsKIt2MGqL7Lwn/uk4yYg6vDMum5lOuKMKJDd4BFDaJnzrby8PZz/ID8ozsani4irTCk11uP
rM9rW0ZHA5Ip1o+eYvi98N665pbRdCS/YaaOENE92y0AEpNirhKgtVl2YI4LWQSK/SyuGDuYLlhk
W2C+XdnbW3SA3NBPGMKVA/fxIoGB3J7wSSPX3EGyC/mubODQBWI5S4TQm+lm6KvSyCe7CEGKUZTm
6R5YIwNP4hUh2XGChvri4I2LZP8J0E85en4coyEQaq9qSkptM30csM+iZnrEECsE/6mlu/gr7Sje
wRpZ0t6Xhc+mJriwn/9j8K8eN+PMTxv4sdfFp1qk+WSUH4g4ukVBqGdqpsWtiYNZ//CUSKWAcKM5
6CGn3bwOrAuSRai7Tba0r590SMcliE/yZiIdcfV+h7M8cXAcLcNyLhb3XByV7sxnhk18i/k5od11
pFzYk7BbCdS0f8dCQGvpbmz81ppZThShshenkqOgR1jP/n0c94/nNCSKEgG+onOikKAdR1HWLdiK
A5vTrCDzQp8naR+tNn72O8w+RQ5sAQEVxbbTE/ROekx2gfdz1FycxbWs2EHekDpCHL9i/yHRSMd9
p6u7xj7GE072FGP+ZAADWrL6g1Q8y69jArOtWWZhqoRgtD/X2dxz1wOPvFH75g8MIza24wdLu7ou
5Dk7dNMa3eu9QIdSPUARPp7BaXx/eECnjols84LrZbfGC5PivBMTtqXFPqh5jedxVxP2WilDbAiQ
/YRm0QphcXnRGBteb9Z+Vxw/oi1DMmHYMHnGP7OkTsXJMslm9n4n24dJWU9iBEcHsWO2Y4Io4r27
QLY/r/pbnRqxIdTXf/gYT6CwJ2E68rV4kDeXE1DqqUz52LiXrIGXBvkmGBd7csHClM1RXGJ9nkCl
0G7W/QyxYyb8yuhJWeg8kAqwGqz+vqSF33o1TTFnNCEXvmB2PL6QWMRasQv6samGvmoc9hXCeAJ4
J1m26l4UQXZDGX8wziMPoHZ6D3+C7DWuuA7X8KnTwLt7jU0knPFME2fl15eNpzNfQOCP0h4A7eKM
glicjc/n5l5K/1nHIiWVVEzfCb40tuKM4RSvtV57oD+4T8DG0d6AHdrAIsLMJzJSchZSkM9QIGiu
6dc7MGILDYygEHtiDA4cdHsK8Kx+WLUtHNBXqDNqlyX0lV/o31rG1uIWnlNxSUEHjlSaSbhZ8lOw
kRVliiW5I2dE00L+Y82LnHi+QwJbTvBKYI64j8Sfg6N5VZrPnhRYXjt7PhG1GQxOJfb2ybKGx+0V
TCrYIq9Yl4cleEbWK5UVbmavaC2krJd8X8y2SuFCmEy5T+DDCNRd/ONfhOn+/3LAjmsjcAmor1fd
5077+F4/zrUv40AyPx1SITYEaBysiG8aXGhTsW3n347O41jXFHnLIhTdpgpkPOS2JC3S3764DRUz
39ymRE3CMaObNIMIT8JGQvahhNU1GvLnZ4e+An0ciYjdeGUZnDyEBfGhcxIvOTurYzay1QZCdeqT
LMTjnTB/38gm7ORBHepRFQn3EpGRmsLAyZdzRQGEIqONCKbYnFr9vYEL2n/hmgMUQ1DoJrVrR6j8
hAVLFNqSj4hK6pqYBRiJsicYLuha8KnAM0Y8dC41JReegysMli8/5NhqFxg3Os0ioZuPQdhL4w0a
e2B1Jby9IaJA3BuQyW0ofEgHk2qwKKPfa6uR2Os736xjINWtkOcfcPFsrymmK90a7IgKdorSy6a6
fZiim036ZQ+5lbP9V6AjDimB1GMBRznSUKO565AMFqjS5v9VFUkOYGWTiU6BvT8zXNTNEen0RIYH
aXG5HYUZYly2LtbJb3pisXYtrB17DBLSh5gIjuCUsuQFAqg5GXh4ZO7u7D3JkmIJyt1/x+f72l83
iMiwilkWjTa/7RF/6er9h2n1iJ52PcqEUXlVnTXiay1eozd57sndD3ua8o0wYYf05UFL1Bv2lhrX
0GQxZiHnzAecuvVbc1JhSw7MunntidoTUGFx3Q/2jE2xrbKwE93LgvYc+zrdfIjXk0MiT7Gf6fc2
gSnIZLqyUqkTo7E5F5V97SKXGirt0tkudobCY7ODInqLoqAfZ78bIsjB9MiUpOO1FqLEJ8913RQu
ohtjCDoZMag71BI7prP/kmIYF24Nxg0E1rpZv3kjJZxAkFkOVECtkOl9Fk2zo13iePN842NIbSnv
l7IekYP6UiGmaIZrX8rDGWaqNHx7NbxjUNlvlGpHHEo9g2U8OuFJfRnrKVyKhN5IJe+DXV3hJPpm
tFOQ/X+USh4RqbRpdFSE29K6Imcj1Zb9d9xD9QKbRuqiPuzNhk4t69DxSGjJ85PCzmF82cGUlPtS
nZgW9Y1Tzvh012Z48exhSz7+vh1n3aw/vj+cAcBYFSjsfXRldovLEjucGqOnuj6S1oZpkJvWPepp
/JapAlIs/axOgivQOZUd1swHbhP2SP9J0XhCaN99r9AIHPrMeY3rguSDSTpuHJ2X2vjm27jgwJSt
Ej7IiMg8iKIJsJXQF9ea3QBdAVNOd0NdR6c36ZYVNKhHTbXLqChbhwY/3jy8cvdGepCIqSXCZ7EP
oMIyhzXnyfuz6EmtjRqVNFIM7+jrHEreahV0HQ3nyTWAaz6Ovazz2sjQjGrJTJ82t/TtjBYhwxUM
P5A/En6CV7EP9+WOTVccp/eBH5EsoWg4rLr9aNaFEbyzd02iNqsCyVIpwJyU/XUYtUcfUNIKHYv3
xxOAZ+0GXDffGPqTEOwrvhKS3VPjL3rghGuVr3/vRXjMqIUrJo/RvK8IpxAdshMitniQr7D9QoVC
TpSyIMbHABlATGSoK1lyQa8sIcAB0YgD8QFUFkxGAOCw0sM38u0GgOG97bDVY2Qu2yjNn39f8QR9
RGlmvNrUqzLcXEvksyTZeQ069Ur8MbyMJ1t8rr/sP2r88zQCB4ldJOrfWHvsxFmyHpxNXXB+DhuN
aZ2N9Xp/OB0dbyoqSKGuKcOFXEIme1dGh32tGMqUAv/i6mJFgtppEhC2Xtjh0BUlrvGPc9V2j3ir
UPQ/5XIE/y7/qxWV4L6w6/BWPdE/QvHILpdxAqFfNt1DlS9qeWhEoUEvbdYEs0mFSLlNP8hBFywa
KRXkJKgAKin9lNY35EBJ28AalnE0Zi14Z3ee5e3mLu+ysR2jRtbqKjOSSLyOOPDpFrP67VSfnnbV
veYrQjt04Ywo0g/M4YFgiqSWIZNHWP05Fz/ffhWfusMi7fjx7cJCM6mQDsJ6Iwbnk9rrj7DaurDP
JTWdghFKipIq9yAv5d00ROsaCVOKHQQFmzjpDVlDAGbjVXs310eUeWRRFJ6AbaQgy540A4UzKGU8
3Pj+pzlOJ1v1fVGoW7t+KTQonMAeFzceVqXE2SST92eDm3Bb7gySGvR/88qc17PqhruJw7Qz1XwN
OXsx0gC3gwcSWtch++XQe9534SkY8Pvlv/UZWYZD8pmbzE8E7NLYzmJ231l7/QSUBtSWtgcTXZbP
SDDiKfmrmzSC9OvOFUt1RDgPqcT9+OGWt8cZ8ocnJUEYQSdiYYRtXfOzv8ll8gpnWx6V2h79WO1/
G1qkWPwqW0zJ0x+/FudlHMviuG7FT1Is6r015R8S/q443VsCrGU2565wSnXM8EEtTU/ioT0lMBfS
XYlJMssZZpqCzDsNdTo8Qzqf22rYoX9qbTlGFq6mHvKHkNTqz/Uuxr910jiVDe8m2L1eWG0mtJZy
5NHwuF5pfIXAGKNruUJ7w4Ya7bGb+JynTmCKzBmsKqZcAtV2Yftkg3I4e+PBZS2xkDDhPWWSG+Da
ZTRMQDojN+d0+xIwXU4TRFim1fb7g26Q0GymGpcC7PVvWnl6XaP8GFBtzx3dsga1DEtiEsSSSC4l
JBA8qAGWywW4l/hy0c/Ylabor5CcxV067aHRI0cx2zoFTFCrJ/0UWcZkp/3zpudGw46bVCHkffHd
qTAq15G+e02dT4w+u7BYa/wgV8u+HSSwZ3WbWKocM72ynoYa3q/q8edm+Bk3iwav7qmj7VcuaMgc
YPuD0SxZmQ/2jtGPU2H/2MKUOUVUR9H5Ixm56Mt6+Ilk0fRkcWYKRZ/zPHbRFcnJfa+qZxjdiq9c
1PSCwN085W2qI/84UV9SVPUeS9HpBEF9TEm2+SHEcfLICOX1KOqEnRky9cY2AoYlKtk6Nph6n4CM
QodQWnKOzz9weO/fq3lO/bYsrOCnH4o+LX/fZFFQ67FR5TxC+uYPnvIhFep5WAaZNUqEETsFr50M
eSXT1TZ5tQS6LobV8gBwWzLgvdFNwwK5ifO4F7jK41DfhuwWHMCFLpW2CRdjtxXtudiPaFYllM70
MyISkveq7A9NDl/DUWX36LZM1mFFm+NbD65eaJ1dl4Uvn8wbdtd1vU24rLWM89/MNMf1nL6NzIpH
vmZ0UgjeCS4HG4mj39PgObOdcbLvjCQbBYUgn5itILQRAKpSLULiaQg/EuDjNee9F4oe+z8NgPJ9
QL1rZijpJSuUHUHfgTOppS0uyC9+ovj+GwZs0M3Heco0VHC3VOzzzQ09qoMtKJtKgtVoqTtiPL5L
ttUqlMqI5yV0csqzgBPuCTBp9Rf0vLXkuwfHaKv6SfXQf0+h4dhv0dnyiDx+7QJJUtdr9nNpiWOV
/pn553TXIohfV5uO54eZ2CxuDITMKLgI66soVMcSGUxnwxnSgQYpT2ZwqBvPQcgT7yNlA/uzwh1Q
s16wQrpMa2Qx0phO4LAsGILXDo4ecfyD07ditjL1PqFlOZSmj/VSnUScZGHvJpUBxlV1Tfe5weFF
+feah5nxP9HAhA96RbhHuRNJDALfTfxMsD7hAJB56AFptAQA5nBd47dALpJnZBW4jsULhIJIp7pC
gPm5rzJpsENCjhogNTAlb3Gd/lsjJoDffxosVt1d7K1efG7ISVTVQ4NBDvzPsKvdMth9lA8xkGCj
W9n8CM3eg31WvtMslvCYLtK5VkDs/IdqHOD7OsShOrcrN9k75nW+goBG9JUKUTPZx/yw26i9KuEk
N3ebXH8rBF0yaYuwkd5+lmV1hsUQ2MqsIMGGmgOpZR3Bh5h/DlzY5KewYgKoM0Ir2nX49+CJy2pe
cjurw6Nld3T3RYMljjwaA16A8bGnUjX2MRzT5y6z4xICFCQwh9iqHdcNWm94Ti9d4+k0PG+HyNt/
RvP1cZu+YCyLzMR9VrY31KKCqQAFHx6HSFXKdZv2wvlTCV5k7DzmrB+MwQYTMtEGmldb4V1lEi/J
YTBG8lz70HGN2rm5He50+ma8XaX8VB35a+JyZT3mOGStUpypNCQIjB3uR78yBMAO0xfWwqrjKwBj
nePZRpV94vjef0k9q5HjXYrqyXFoxLgEzleU5v/3Q9PbBvyNLHjLVP4M3P9YPszE5DOXiN7dbqss
z4nwFwdmDAnDotFu3zNpPhzwsxFLItjl5CxVMQ1OM5jt1p3FnSHwLayI01YLUJ7zKAysydf9qza7
wZz6uwiWuB2H/a7os0r673Yr+3jJsneUymMyIBXGkXq2Y34KiC1IpVDsJRyQusP7tpQAgZ6/8lEo
RE15w2uOIZZ/ZQ6Brqfj8mOoYvi/qNvvOgQrHbeR+hVLRiAK05f9jFp3XS/+iYIigumoZ5zcSr4H
s+ONOHg3fEB9wwEZ0qNA3VOXjzgiqJ3Q05ssGHWMNh+nAz/V1OkisroI6ll7r3CyftFHmVdKjcNA
X4AuBh0iaec+rezgOMd/8hPHhYI8GbaRbc/gBfD5ZwuwQjnxp4zQgE3P6/4EjC08YvX63G54HZqq
LFSqZ3Cb0Lv7RnwqlK9DFUZkObtseYcd239pKNwjyj9+QL8SJRsJVUnMVw2GxMeyeOZklXwMlW9Z
Ljs=
`pragma protect end_protected
