// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qaZEEd43mue5V3S11nIgdVY8UTehCzONGbP7XBa5bhFyN/6nXJKWMZGA2LKCyzje
tFK6GlsYgi+C+xbLgarrVGuxP7paojoglOphFFV5kKpP/VSERg/mq1cXeayoGx0r
RQn/cpKfxYDYUOSYKFkZ7Ef3LldRrLHfuoYPXeT37dA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
o9FfQeq53rc8j+eMJLlWz9v1O7+Svbhg2cisz8+XLYUti0GQphOncSOUYTyrdrXG
0cMgKhyI1e4ji8mytNg4Y2/xXA4lSl29EAhItx6OPPXc/ll/RWA1HRSkvBVu/TrN
oZO7752DqUwx8NZFasI6AcrZNXPwf6CjS818HR2lncwVmRtvevqz5+7+p0kxxGWl
oNnlJScbP29EWSThMttcgG7cYwgNE//lNpU/TeHbt+sAQfgWucIq8FDi4L6YYITd
1rceSmoABfcFL9WGIVD+G4H9dJ2mc6fosFDj1LYSUqDSAyd34Lb6wMstls78GQjS
oEeNloGX1ndHQjlF2Hj6p1bRQbxMWdUObH6TcUFIkrB+Zx6oxuhoQ7U2qpvS5gSb
iaDWNHzCE2V3HVcphr38r9IGkxa7FiyQHYxEnggTFdEXcROWYsaAQx2RegeVwhxt
KH4CorBbFthTbP4ZFu+lwX7xjdst3QWqukqWMaAX4YiDtsGUucb6zK9fjLCTY2ma
Ck4eCqfap6/vWHOEsA6Zuax9aFhaSCQ0mrxZHJWgtznPjcUpvSscQjGfOva+SzFi
jd122QbdOMzOONVhwU2lR2V9bRV3oYVXhKs2jQw1mEaM8cUxAecq+78mvXIgGOD6
yZsWBMVIrP4p0kpArPjRMPVt/Q+4BZdYlvwi0SBr8xJ1nvCbTsUidGYY1+FV8/Kl
JyYnQIQG6mPUAZD3l7vD56+3Y132sf2ybVhVza03w3iNM9/AsZCWc3YXYkEH5bGd
IUOTekhtXD+0gqn1VPmoOg45uay71WjjXeut8hSy41VKqDhk58aUr1rxMHR0ieZa
Dg6W7BlemhCFLRTUZp0B1f0SXKhKnTySrwOhiQxHvSi/PIC665sK4T+Spsy2yZlR
PXdOQeV08UDUK8IAqQwJYMLfaQoIU+AnkOxlOJ8BYzkB7/e3P6sJ8ZZ7jNHzgK1g
/2mzRnCSb/U8urodcDz8Y0g9irjFJ6OY/TJf5X5UNVA7YgKJ4WzjSYuVvibCSF9a
DYgLdAyKOuMJgwI7pptYy69uwAga56UxpIPH9eupsLxdyQnvwXhq015RN8w4ITQ2
6RQ02f7RWlPQYB4KY7/QEn58dGJpdEp1bqfxbr8RN/hp3ah/UUEL3Qf7pe6kvhID
VUJeygkMF8wV9B0BnUKgbVw6PZmZ+hXq3QxNgr91XbjF8X1GvKYKcdnGShX8CZpU
wWRXCB7YZgylNiKuALHMVznc2yZBW73xBU/ee8sqxMfjNeDKgRThhCnoIT+anBOV
Wu2AfhwEvd+QmhVfxZhKcKMthm7oJnQLIMUK075a4KZStjLMuUxF5hnqOuxclZW1
Z3h1nlB7m1XPPMM6YFgHDPkHhPeSM830PVvN3HYfzK31ht4vizm7BdclsO5XMO1Z
XTkWI0W7PzzhcXEPFeD+3n6yHjKmMpE2VX5B80p9cUE4JABFDRyAOwfPgzdoPI2J
89PhWIpmCVwzAlVRjHkT3X8bOp7takA/3+vYFcJNisHVDTyrq2uD3QeQ4rXic0+L
7Gmitxm/JeB8NmCbn3X18OOCNOzFmWkHw2MvX5oIlkQgJdMdgMlmRhBokscJClke
PrmM4Jd1vsyY7SgQjA1ix+9kMu/17HUl86vyFPcUoo2MdmOSIZYtrhE6K9+TKfVW
oI+PaM05hctWK0bt8A5iPDuOAitB/VRNu8WYQjN4VqXtijgT3cHe0nZef6q1tkR4
JZE/OcvsxObXqfYWOVb5NE6J9zYDumkdeP3Vjp6glyQAUK68F1oE+k1VxZe/9GQy
sFxMEyLSIKRQJEEc/6qDchIdz/sTPiZak8BcV+H3KZMTyPNzKOMCLquLo1Uk4ScV
NpcD7YCz+KhsPyBdt/ISPmE62w59ApntPp1pAEqjYuED15paYdgxpwxy7wfFNORO
aBMMS+PUh4+BZA+pNYsHtKnNVLfYeN0TWDkXe8OYPKjyeLxn/fPcnCz34xH9vmWr
B3w21ew8L9aKxC5Amt3bo1rattQfoB6FV1nuIWTRj7hqM+/QVboWgJQYxO565Pos
a3gm/v75J3M1Pqcu9tfYH+q5j9029Jy8OsfDZ1wZuX+PeKnUMTvymR12hF7TQY39
2M+6ipGp9ljWJuGEnvhfc5VFGbP+XrmS+M53l3Cu/5JDneBW/ubKpijLJblFrK19
bLRhyp5LgkSNM2WqBgFQhAl/klaZ1eu12FNUkJ+jenAGVC0+xwBv7PR3tGJ8sSQ0
0zFsvYUt624cnJCnZggWQiPP/UHlpfy0sbtRPRIYMe7M+IOTgqX2xpySan74ICHV
dQvBZIObBLkjw0ZhpfvWSKOebVrPxojR2+SzS9pKPl3dRN1tOcRX7qzqUIRF2Z0c
iX9Bl2snG2oaiN+UiVKmCB5F9lLV6KDlrGiqXOLmsgQyWDsqmCazyJ0GjNfhxshj
mmDf3u8SNzp3NJK29NCUdxpKdWZR0vSQ2Dl4YLQ9kQHqT5ZDO7IFsz6krAyVeWDJ
Hl7vLdQpXKaAA3Gm+sxxrN7Z0kcYOlFM1MCc4kqFSCamGirm6uNxyp0FPj+f1ADC
kFAxnlhBmJoVvHPq1ihHEy5xfHaOjTHdHR7o3q/Nqm1HvfyBK/0IjWN/87HDCUti
9aHke/+ZKoC0iWEAJAylS3AyxMhlGw2NoMzoI9OStb9grc0q8kTY4gmz2jnqO0WQ
Qf9haUKdL5O7LaraTNgDczPJ26NDIdv2VZad+jXCBmx3sdqlYHBpPjm/kDHfCHZv
Jxhjyv2AcKIJ/gn6cTfUwZ81+IdmSI6l2qWCLyVAX93W7MM8Mjs/Io8Q3HvfD8LS
tTh7yO6frtk7Etk2IwRGyFGiCqBCYzsfaUOsJ+snQ3CnIH+DzNKKwXvkUfCP3pmx
s9vVrnqXAyHmx8PBJNQb4tE11s6S/xHV+HAgDdb/XCr5+ZLJIiyxvY4xfQqqspuP
QNaVnGsjqekI2NrhtYLMQ9BR78CMOlY1iFZvs5srB5YV2uChurz+Ly11QPVF6D/L
0EFXFCxOM9NCm1HSrFGT36LIRnBzZEJXIAbtEhYMvwmBdLykbgo2XJgzovI1Lupc
4FWsjK4oTFVMVLa9Be+GA9GcU5ENtP/jxy2LBsMwa97mA2WsZWPfcvorz9mgtLlN
QS3eVhY0Ske4XoXmooQOghZMhAdPtuDO/y3Rw3hWQ42K4JrhX06IKTlrayvQHR6t
0ocW6kqZsSNFAHm4HP3Hz8QKqwyuKTKjdFaDIzTRLLVHwXW0X644ZY4RlKV3+hVX
4MSdsqufrlNiCxRNXgCnETL7Lsj+jrMoZTbt4HU5kK/oblFLkud357t4gD289I0c
o0ItzeUlpy3hxTg/3NjpKKjZG1ez54yxLypP7xxVzPPlfhIKsDhHsoFMUAaNcwg8
pFPV9+Rs99v3goF71yyx9CbqZ1d09hC1k4ysrLRIMH0MhwwI5bb42ZzLnTUvTuNV
wXAFrYGpKD7VdScKPNAYify8cuDQWrZogwdODsfPJkxbCyFkRivyRVO9KqbOkRy2
Md7r2FLo3wBmWSMCLGo3VC1bCtlrU+Ci+48Pil+nVotGaMrEQ6xFonwKHPEqfc2w
jUeh6B76cfOuRToUs6Yjf3JM36qOIftZikpIU5zfrfq3pNsfyAM+PXIy9aStpdQv
QV/u6mX9Ow2stFmaMTsIJkDj1yYraEkk+KesC3QuBb5ukic/xbJpcjz2QyjddS67
cvanrjlx9ViDj48YzOFlV9CMCovvuM2+ZA9qSwpfxQVtGZGX9NUPE8IRL7macZuD
qMzzKAo5i60eFgSPNCFvu4ztk/gyYox+YcwwiGB0i7U6EZCZhhnOgR3PtlAHI9G3
zlNu5g2mRYqddk03TyInlSwX1fr1nytenaYHzngA5aQ9deXjsYMRZnlVeCYSjwcm
qb6B0MoXLiQ93xDTPAoljs4QAfkHjWMKaHbDZTKuRN0/9XUoqEE3g3WEC8whpvXt
SQi1e8BbiKM2Y+/h6+iF+glyMEi+u+XuNhzldI4StxKdL0dtrgRBzmVIjRT3SpbX
rFllwiX/G9Dr6CwdNU9MfJ8hwHHKIn3CudKZTUgSKt7xIxQ/N25tMW5GzSxfrx2X
cDUzIxP2fUVBGtS52r3a0rRZw0QmeCKho93hoY5a2xA=
`pragma protect end_protected
