// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Res1Eeayl85T4qkKZo0fvGF4UOVV54dXu14mWzCvw6cwkGmZkiVGJapDTG+ocLE7Skm/twdQ9b6M
GwevrNZCbGDT9PwzblnF4In1ZK/MsGm62vHw7KGNoMnw7zYs9h+G35BbbMH2f14/FSmx6h35JPuG
k5QwC3IM3xIlW52Qoily1ASYHmoHHoeTYgKRt2TlMlReaJbYE9zHszq+LvLVXCLXcHqFMq6f6RLj
lrhvJeLAoEdFfwv2d1mhpEpIkNLgjun4+D/P7deNW/f61LLKk2C8hSa/iN6wrp9NWuhZBvvrtWEn
BIQE9mwoC4FlvxB1HkFHQGsAcQ1a/JSQjii63A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
5z814Dpzg3EvxM9UBp8xZ/r1wJ6pN1FyG3iG4Yjmd+3zMqSnCtxBHbmw79M87BZMlkC4xD0N9NID
JpxFDJAv82gigmKBQPIHeccfMAf5qCeTDNfLSqy2KBKXuS0AhXd3cE7JaQtV+KJm8IB/5FAqnIeU
B/Vev1GZJV+BfgYHLi1cLmTHVlE75D5UQlCT/nEzGj0YSkOY9FmbmihpfaxoQgg6EouWZ/SX6SE4
wIAcgWD/2fTfMtYkQ6NMneoWCwy0z8zd8CzySCKv9FKAv0qqCPO0x5ful6gENcPxff6u+wdTFfaH
SPgelwkPfVsiujZqxErnZ4IebgLzbmwySb/U6mNRQ9nBdJkwdIkLD+CiAMAoTH9c3WxQU1v8p5G6
GOdnKnzuwbxByV3AJkiwMlMnBMo2n5WEbQnvCACa8SX+CYZ9N0bFaAErdSV1ZlkTRPqd9K7bWPBI
WK6glbZnzeu7mTXjbxCT3OR8hMSHAasxJGjaHavsXR9EedNuSq41gHV+ZcV2CHjXCtqiGYaD4ykJ
PECc4MTUdZiZqxLuLivRm3jkyv+8Cx+hgbHQ3nqMHL8OJupvOtXwTNrHS+jeCPZur582v8KqxIAv
sQmn8RPF821YeDM0KLR6ez67UYS9pttCdJjRVv1dQ8gi50s+5u7Lj2Sl0Vlw2IroOOt49f2AAzuF
AHCSBeW0kR0C7cwaU1C1yqHrfSikPurCqnWpiW4L+oQnbj9rovuWWK3G+YDC3aVd6XMHd071HRif
kFS7KK0WdaFGOdvk0LYO5MM0d29AAcBYSQz3egGFYYAtWCADTAHwW4Qb/mhW6T3VECB/eOUlQblr
OuN1sHnHTVw9VJLhj2Qh4TRpzuHotOq0Ov9O96O/8mEDqTZOPtwSJxZaoKtRpzP7PGGwlnSomKin
/A9kkG8Ee1Y18msjynq/imowW6dJ7G5J4evuWURtw2SBOHFKOoZzUcfgPnYixnFTIX1iBkmbhtn6
IwPAzRd+XNAmKIAoEWNDZa2Iw6jGKb3DPFKedPbtD3PIcpYA/00naLv7kpdDhAbgrszLUCPh0P4N
q9iQ9k2Y6eYE+/Npch03nVfsuT/UzguRcMZ9A6QdyloF9+GqkdSqYFw/MN0ISXSpVNM0DDGu3/dc
9N5As9akdBtzh6Ba90q+3kscFf7208dg67rEn+yhF+N17DLpVKeje6yIaGKskA/GaJaYRby3/NyJ
dCgaov+OOqCLbpPnU8OyzHvqCxrbDv+Sfyj/0lpxGZmoxblYfz9FR7/vlWJj96Ld/hWXmiTr6ygX
vEnEExGKMgM7qcUhACr7l/z2B0YRB7mtdllaFfpmWYSMxWeSJ1IQsCPBwBw4jeNxtyOib2WLNoO5
xmmiKM3TiS9MfMZqaFb+sgou0IhSlwW/6e0Qd7CfNXFVOS/LlnOwI0Z1qAqSiLpGxTIoH/0YeWWj
ty9s6IlXL/2wlwW13DaiiyEPd+jog5jT/e/EUZSmtbtckdhBw5/hYY7GIUDt4v02rtRNVZX2bKkw
C/c9ETk+Z/LwJcHeJvkpRJP9LLbyb+NeMHYT6gKSBvu1jQqZJdq4tOG5K7iI6voZfMT62ooP5RNX
pJCAKU0XlA03XIEVXWU1UDv0YSAhItn9rdDqK/K340LUXkqcPuxk179IWXs/T4e/2DI9RuUOiaCI
wdI8yvNHajgHdSPRweHcL8P0VkIpSsC9HlHq5WRvD9tkvU1jZUi6MElY9M1gYmKydl722ht+aOxD
CoG987zBKUI8Nkg9gPoGoQOoyVV9E0C9Hevk9EZBMbnUbYgxqN3L76hUu1eTTNmxfUNNqbALLU+L
au2aTUvDy7lCIAtp3CkFR2ItvtXhYdElZCJOfRDuBx0loi7Lq5gXJZyIjMeTdnZrKe6pbV0kQeS8
1bKgHH1nWvxcep1+2ZPFpmn6D4cb3dj4KXcdNi6cOMQlF9JNDO17EedKE6RKwj4a5csi1+gMDIz4
jRDZd+fo1LdOyztmu/ceWyeVPN78f0Rwj9HveFxywAsP5cx8/OpZ85DCUhYt7Gdxexk73gdoFeRM
eJwj4KjcXXXUW3P9qg0S1PHF446cD9KlM3ft9/cLx3vFiOvXeX0Y1bJc+SHXWmjC95kY3Ok0t6UA
Wwqw6LJkf7RYV4fN0ALQDL6q+75/qbAM8lVLCebhqKcVv4XHDiQrV1SqgaYkT01N7dpw7RhvR9nm
NopHqVf40rdZXpFCApC2OFP6oCbljVx84dUF2FBR9dLHY9dt9V1VLBYvJCLhRp5cp1+J97d8EhzN
tjA+J/gag7pKCoRCQFii/t8bRNWwilCuUFXRkZu4Jv3zW7vQtgNE2ax4RlMGFmUMcfQB5cU/fQbv
pxUKBPpvl4CPe+Vr4nEAoZhJVOI1DYeyIJQBG/OjsTjpZAnzEPvc/zSrhFo5KkFz8lCLbqzU7InP
Nw4WHuHwm36q92sw1UNxcBl7n31GCobqhYSJief+dmwZkZXadh7f4zpd9/2qUKwTt99SKz5Ic0ce
vg9aaUGh+IHpyuAsMPbuMv6p4zKahP8aD0dyQa9nj+ewu/5HjhLMzEjIxUXwEZF5vesuv9w1KHeu
IPXYsGi8zKOjSBQYqds3pUZg2M5oyqEquTTNNuGwgAaLHTROo5WWXcKwjjDlXA==
`pragma protect end_protected
