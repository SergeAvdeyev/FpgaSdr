// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WtMiY6PNSi0sd4al7NHzEt9LfrU9dPTtJ6NLpZqe+GJKdrgW0Z2BdWmduvkW8Ipv4nLp7LtzTmZW
PFt0Amcy5aBuQym8XPKk+PLUw9cPsfFkPTHWKQgh5yYSV40YchrlDWs7H7SePFMKyoKDY7urePnj
FrYu6Sr9JzDMf5yDSzX44T7m676NuWjatVjr7vvkSF5fIYxLDSdEEU+jJ31Uz9Er7iCOVc0OB779
4dzCHPcqQvEC8JbstEVy5kR52VaOiUaofiwix9PhH8J6C8z/YfHF4p+iFT729DtltV8l2+zefEqV
cowKfd8nx46fN81dUSLXUKOeNpVqzFtzPmN5KQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
MTIE56fqtCVMlBIE43f4ZqYB2Dn5PTBtQSWagv7IJD8q9FPPAG7rN2pEkNfv3xtqiJI45o4JFIdo
QF6l6EOZ2mObq0qTT3jajlO9zm1kRFrOmyDIYfJ2f2/jGMYBB4yymMJ6eNTYHlotO7L6b4VMZYUi
sFLNq5ycmpCqRTLLRCi/6B9aLwtdm80sdotvF/CoyNcQiu+ol9/JnZyyHdO7ED+OpXOQ7Ig6afrx
9Jxb6bjiXQ+fwxtpNt/yHTDiVmjPRhXyC60HCZ+/HQrJnt8bTvcdKW6Y7URfa2tVI5AlPC/5qQAZ
k2kv4hW29uEnJgjejiWdiTu0PIlezJlObzCm/nBPbBKzsefZv/EyEvIOfJjlecnS3POlFg6mCLJB
I1mLLLY2xAgNCMOMBH5HoEIKS2fM79K6wlzIeVjIfiN+KnjgvyW4neHiq47bs8x7v5hT1VlM5Ren
Z2n7srxMBSHH2EUTHCYRzTaqHEUWTjZvl07U5n6VCv1P2/StnLPVz1MYM5WHg1B05kX0bAUk5BxB
Rj0sqD3d22YrZE9Ecq00nkZTiD2j2jcK5mrkKT85R1CZv5LK4X6biW1leTRh/GFTz4ke8P42U/Dv
hJFXO++Fsy1VGVXuT2MguycN1wwSD112dBxV1M9pUbpRYKFjXXdLX9XuNZbSx+6boB8M2LRx3+IB
pmmQOdEZ0wuE8Xiveu0QZVjL1bTqmedUPWjfj/hjeZGbKengzFCEf0fiGZIjyhyCSAIsTuZInW0e
w9wZQVoiu3QZtUutvlqhGCbqmyQxNDMUffru5NsEBamIPOEBeJMJZnZAt5rKXcmKlDpSGNHkUhp+
TnJ44xWXbmSiXElq8vOd0jYHDtfVcnJQ4rKQtVXafSIXiQO97ELNUH0+djvIL7Z1sEgLLf8v5iPk
PAU5UKRsNq48SxW1qVUSep5FG7aqWx/2oF+vKBxOjf6zBcLW4I0XzWmfGqObRAu3sd1aOFPZge1f
YVIb0diPdl+NV0C1DhFyChY4TpwAxZoPUReOW5loUz3MKeykDNWQhFcGRcOxlaZ567vxmcvbB7sy
5sq6HMb0zKAxSfGpvsF9h7huPTsQzHnjq0aemeC9HTpgcqXacKWwm09FdNVCa+fj9dudPGEsdMTP
Q9F4Klp0O128UMTtjLKg2Y+olG/DL1cuU5FfQssxBHNX26hgPRH7fWGlbDdeCkFHqNia6VP3++i+
Ixy1alWtPlFdctghCTJBVjVyplOmtDQ1EXl7WiGji9/mgQ/Ym3Gq1pBoq9pajInnepODcdXDrMel
tCAQC0ZL6wifxhmWpnBzhHtYZzz8n4b2tdeokY6+wuHHQhwX2tQH1HEC3yfTxBGJEs+22bvFVfJJ
1caQb0ZG2Ao83nnB6ff3jWda1oZUdUBU/f4FuhKUOxP32YfLfM4Jc2ZxdlEsP1AC2UBLCSrr+I8n
xSkdI1CPiRiYhO99Rk35oScQzhRNd3IR1Y/7oWjVvsGxykpXwvsziVsQfQCPIfrhllHfZz9Cgv4l
DPOpX3JBpByDmijMqUAG9YR7ps6rA75AS05a09DVUZk/NlGKnTGuW4REXV5gdaJdC4rpYF4V4LLI
HWRlJBVMXHP4hfXK4+aQG8QmIfqFkXBZ4WBcfqAeqSzhmGEKhqUxfV1W/GU7q9WdwWmPoeAraBHr
0n3/rfBaY1l+HUmHkoNcprLs1FgNAip782STkC22sLsJnPyIXGd8OHqNlKediv+bDvjPMIxUoS9g
yWbch0uVRGvU0H275h7dbWLeUTi+1LKoc6tBb+MBsPH2DlMwbA+zA822EHXVvnZTjDtFgSZuMxg+
hh3iLmXkRE7ez1/siLthklokIHJNBgg2fyUZibAsioTQkrOQf7KvODWAWQfTNiotYWbgJ9qi2FTH
Pw6HiocHfmkKb7mvjt0+MEDOLAaCvckhosPqTq3P51MfDaDZ8NJeegrUal+SX5RCBVVNkoCwzQa4
JE8QBADj/382IabZimrWz+hrXPwAjWw9j/wGXFwlXo9kUsxH0a/0X5ByeyF+DM3akrZPie+Pr0iA
dUvw0NL1f0qu5xD/l20HhzAReW1qiRNgsTLxQEurLwgstKOE6s8FRz8Q3pMaEGb2tP9bvyR66OCw
3fD6kHbiaho8bIH745BQZwglA1kJ9MGVXS9ilFwajfkInLHDsfOfpBCrjn/0eKItnyq7X2i200uz
yw8psgRsTW46fyB9jagMZg5WeE/4I51olyBD4SKmr/7q4yW5h0HbWlkTjc+nm5Ifj8qG+GQexjIi
YcbQdwJUWNeHGjj4vS2F+6f0x73z1HiRks/QA4e3gMi9qojHX2xbEi8t5OjY9vrV8c0Xt4f02CbB
iH/JZOZfH4xQJtQ1PSgdpRIRedYmHuLfOMTCTgwfA7FbgL/TsVGdjmCMLn0+l17y8ZfZKUFcwWiX
qONJLW+lCyiR89UmaKrClDmFqf2ghfXF8bfcAfZwdI22BdVPiny2UpxFN40VJ3Ccy6ICjNfo4mI0
VSFr7Ri6y9e8I7afnYr49LMB4eWM8klw4TM+rKMWvUCIH6ibdo+NJwJQFU2YHgZHW1DK4NMqX8Xv
fHxKDB9MmHiMrXzS8EKzUVRZJ07+TDeaK5UQq/uEfzG2Mef0XV4SKTtw6fTBnlG67h2V9uYOXwIl
Ub06rbdQkhuNgc6OeHos7ZtnCzPXgtGMqP8uWzxVAMG2A+TdUk2u0/KHdEK82/sMvL/On652ou+v
2WjeHbwqfmtl9dmfHs1NsKk8/TJgsxB7I2nY+M4KSZ3BZr/v0ClvQPUfisZgpDluLrjvuEYJfFKh
9U8AklsyUszsUAeDtWI7HTgVC0+CbsYH6DwiiVVzzVg66Oo5/y77LvtgcQps8fvLQmQ3AoSvXRj3
8wosnh/EKAEseKPPQlI+UVGvhyQH5YoNa3/TGzTiDBoCYWdMOO/iNEeYk7vS8D+A63sp6k1iO4nW
fh4xO1GeUyO/lUfitZYGCCzU3+Q28DYyEVoOAuSchZEcT3dDVhyOJ1yFlkJFlQpIwOzvO369AF6B
ofmtS2uZaMlux+RSaF9HN32TAo+sqqPYkpBryCoVfYCHY0gdncLMxCXrsg2m7L6Z9l5gjUjwC5pM
xH5ruGBXF0sU92PRtfcptgGzH74LzvPB6Fw4V8E7QHwYjpKmTN5KzgPrFmdfhYVTTKByuVQuIuVQ
Sa454gjSJwKkHxpyzVEYB0ep4Qt7UGPtG1jXPOzDx06FINRp6Za/gwafEYUKfe5ZScBF/JYH/YBM
gs/UD1dfRZK9LMxTdxaKhzpe8N6oC4GnOdbpeTxxZ7jRXYl/YYoSv6x83nGEvo8MCXaFf2grP57h
qXIANCSqYdnFUd/YhbVyYl6+P6IicgTDkPB9fgH5ctSc2/HFOBI5iXnzGHtLH9NoDvcYjO6CL06i
hwwZf2AodetrNX7ysKs407n0FrJf3lohFFGNu3HMONJ0KpnPSk4c392fPr9EbglJzvQ8LqSntMDZ
GLxU6JT0p20VHz0nCMxfqDI9OzlLv6Z0kzYMag5Y6/tcMjiwfzbLhMudHZ2RngucQhWLdO2t2OBZ
5TgemOdxKuym3ht1UmEFofs/cE8Xvz5k9buTcpM0GN7J50dOWohwm8IeihBJNcM3C96KLJa/DdOy
ferjcHI3jKFmhb4lTzIul9NPCumIDrn9+dU05usJJHdduv12wGXVTSPPeV316+yLSpqNMivNzkCX
XO0OPwZjso/8qDdno7ZmBcrYtWw8icJtLdVvh8TuM1WlQhtDfhiTQDpIuJ6L5nsYsjcUyffezhrt
7VHZzxCFhkr/FSNpYMMK4NHCrhzuHKE3hx0E08X95PHdC0TqfKHsmPxVcOHYK7GtIdAXmQkeEliY
NbZrYyUew60yRAKyC37cYr/zn4prrUQEl9+a0tW7ZwWXtj4N6isQXs26Z74FnM9+1eX9TslHGzNd
zw2GQw82njGehGD/6uX2WHogdlNuT9ikmn2ZJb+Wpe00Xw35JPK4A8sOzYwrJrIRqowDP7NgvW9j
lSGbKaEK0vTqr7ZYNqx1IkL1TARIb48CjNuSCRqeGvkObEDmdWd2JEcLCw3QfbeTmmrWsB4wttAM
HjGtb6EWSUgl942AlCcgIBXrJHyDP3tcHJVqQopDTbOyS7XG4kLeh1rCRRxImWV69iQwzozHgTnG
DyEk3C2vXSIo52TZb/UKhBQipMv3+ggQUVAm5lpbAj8PhNk2nhg2wem0UI7J4AsSjF1nBXrjS6av
1J49aG8PBdtBvKojD0a/iKeEFvbqMx+JwQmEv/lDM+V6PFBSaMfP2vp43UI55aQRujZ31UsQP+2X
eh7EqNi+QGQl5EkMfnckeyrwhodj2k8nII3nowSNl1/dKh+Po2pC1PYi+iSaItgvHsD9UGDIGLIL
WgFTA8GVLm1knuN6kLwRIuY9lNKIh5eEOdkts2wqxoTGQyQQr+D0U8kttNA/djYfeNMJLoKA8Hgt
GKcsM0RVQieWUIQrFKiE8IKOcrrH9z0oKCuRRMV/MG1+JldQ78BX76Es/hCsXakI1Xk6nOUeZrHg
mHWkoaynB8JejJ6Yrth4WiWT/XJbQYvouLfhjt82spbErJtLNzVaX9AohWCMUlwNhUpIcVeDKbZl
KI9GKPk24xiOU2BTl257kPWqYWb9x0rF/MHgTugdlglUUuxIy1TVWCfEx5ZvEi7+wIRddwgrHEgY
rDtGldhc9Wrn/hmK+F4OVN2o1LY71S/C1lcNw4xjSkHkuU+kDG32TcAECAfwc9Nku+p3nAK7fKqu
xvn8nMpj3x+U9LDaob2OUlDONZwl0JXnkkvP8K2emn5vx+Rp/JVX24C40BkIWf9dQvlYNWdocFpZ
ZYgwk9AK6byy7FQ52P3qe5Ohi51Bl0xYE96Twb2bX4HuwJUyRU5Vppw7b075COlYhx0PJVfXTZnj
EdUXcBio9G8EqosBMsnETqPjJV28t5f/WaeVrXhbyNJ7KzzRgkCoS2AljrU6WlIlKsQ37E4Mf+FN
rJF6rEnAVZilQ6fH6ngvuLSdby/3/EzMPtPqg/po+NQa26+J3f7TlML1XecKs3jEgkyK040YGV53
67fOmSzsV5h7MGSidBEnT+abkM15YyHzxVszMHlbHrobG4svP/INI7thKSeWgdOZaYyGygLFlka2
Zp9iQ0TbUWTAZvkP8DJgRyCNh4o2OA4HiI0NjdzxOgDRdOJxTDLeEqTzfGtym/xP35tSRNT1MLDV
DxpXT9/PaeDtcEzJ/P4YMjgMR7C9nJGUCE+1qOwdyybc/bxpcE1ulD+xsUxxltBC7hEK2gv+nWLE
Y3XkZHxukVgrsXsexlictEoJb/63zxD9S61gkStZo/omDXwTychNKsD/T1LgUdQlz/0FvOyyx3Mu
ZgIs02/zudmeH6UN5BjpRdzdoVnoiXaR13bjBY8c0qKTr3tYhkPMV1mAtWpoWND00xho0AuuzLX1
zFrsQNTlg09iMNlQLuO0eavbKhzcWec7cUSq4INxBMNiMiy001cJ2xdjvz4rSoX0HZC25z/V7Dao
jGFnmub77UA5rwC33hNYKL/oKxyFetaRmvVo7iwBmrGE4n8Vq5YUd6Y+cF0Q8AKRPta7UyEINc/e
RoeS+d80hsWabs6MuZtq9zWXZFiIZznccJkrOiSmLqXXy25Cg3XJhQcjBVfV5w+HqENoZMCSGUm/
OkaAeNXx9/lOulp0toHUK443HKArF9tYj181Pi7slZn2Oa8UXVgyFHApH/71a/Th0pmuCkLvjxHm
Ft4AAMFP0XwNohK24dTtm8TfgALHaLAs76zyoP0S+cqMtOBvYomI7elk5rTcQgGtVmoWRusXbtOU
uUuo4d4mZzReUlMhp0nXSj3zpynuqsC2afkMonKPx/0XxnzT6sECVef6c0ztJ8F93E9SlnD6ugPi
skqBmdt32zTnRnXDcD9bNPzAb1jnw5mwrjJ2Ty+Q/ltvCWx5ckIjAxyeQ5swL3fq8kMs3wsZbkyP
Iz8IbayQW8EenQPllcOgLZXfpem1lkiDV8Z8s0/o/9LZED9MyHN8XAvN/C+x5yiKjBw4ou7yhVpP
vIWI/NnaUN7OR4g+cQp+KcMvijXiOIdDfBjYj8XP5CzNBYNGg/0nJEaW+zBZhcvWoOISl6bvazAe
oihnTfXS0cuD16sGitCBLhHf6gCqrUUI2BFRZpnLqkc4/gZfRA3wcvym6buI6/uysLT3sy9Hjy+b
gVdx7qRyyUUKAZ6ehGKZy5D17QZOW1fmmWnExZQE4Xn76N/bsmX0l2tQgc+Alg4+B2CHg3qyImz3
6do9OxcRHW3iCZixz4TmBNpvTeFUFqrjPgbKw/jRHN8bm267U6aLUNYtcIJXF6PRwRuWDPBWHurv
idk/2fNMkJOThDA275DKSkYeOcCr6Nyr2vTF1PdsOLm4eoqN1LdQH73wpmhns5Im/TKThw4YdRUk
gMw67ydB4aW5zyQVZI5XYUuSDM/SbL2CupH5eoF2LSKUOTV5Dw7Cq66IUIAJGmO3OVBc5gz6B25T
3+/1XE1vUWE5gAXhxTWjP8+XpcS8djq3wPzlDUL2hDqiY8c5oPc6ijTPWrXJDPQKba9pZ7xYUN5s
rOhLB9PWxYM+zEBJp0Wo8ap0aKoLuheVhXxx0BRkSvz1bxt0CKvmhzW5GOK1xogIfyRZ4ZlX19Pk
k7JsckLomkjxsitjkoxzbOhOuaV3eWDRAefHGbZwfXbgHsMcOeIi2XWH5pNTbjThtf0DQhxzYxkB
Kkxg/nCHE4Oi07dlntdSgec+Du+d/GW+YPwTVaePr1sFyBxJDXqpi4Cnk0Ux2YWpGMr7ztqBSlAU
sOOZBYaseH3mPoeko9qbKbtUVd9oKr8FmrYGWnHb9XQG8shyICZSWc1sBux/agDtHRJu6uY9NBYy
nu6S4yh0KQEHs5qFL9ZK0KmvfaGQemUjQXKMmL04V5QioCAYxbUurQGDvHoXzanbhGfL2Rflu0y8
hHIqJfjQ/GpLGXOsJMpVMh+HsWDbnW/XWvs1siUe5DuP9XTy9Oey1K4JluCtOq196TQmJkbsr+ks
sLxXqPhln8gqfMSyghX1cbpFSeJXzthTqIG3LFvtA3tw4/dBp8N5GjKd3+BVSkF/+J2Jj8jfRD32
WGfxrRQnrpKlcCCqFPh/E3KigI3PFDkLdJn/Cs4TWiqMxmBfjHyQMalShcdXhmwF4Q27BKkQ6alO
dEeXcAcw1nHfZy5T6Q9MnQFz2GjxDo5hLFKHhqjCpJSMWNmroRNmg9/QmiCQz6ky7QS2JiwQyWDs
Ot3AOzPOUi7c6cAIeggsoW/U5/RMOfbhjXr3bPndY1kqzNp58tWdZaMbAt/cM7+QJ1Z29N8w5yz8
GSpSayg2a6rvYTbRdDKPXGDvHlvRDtuweW7U+yNxGK2gxv1/7eCLNW0d+LWo5qdDzFaOwGCon/w1
+aIznIlqy+xk4IVd8TH5DY1/BOw1Mt8bPgIvj/i9I0UGIQBAdRi/z2+sdNj7P29JMtzOXcMx2KPC
ASNe5sppRWBoACpqM1Vp+8K9y4ksz0698MV5kd4pacl+MsX/9ow/fzN0VI3AR0UFRiAKc1RgFXAa
oJOIc9WBL+nM1dMIhvfck1k7hGRHd+oeOwy5du5x++XtE2cMlnHkmfgZJuBGObvpK+auU9lj+TRF
IvBrRb9V3EwG1sIVRjY+cRwALHvs2IgrQyMUX8zcT2YoOpS0/Sn4AKbbgDDhjbo/mN53p4jIIxj2
Vb06DTG1EZLDkFSPLa2dVfueUnSDy0zhkwuG6I8qYsrjQZ6TNYY4K6wYJhLjOa9owKlhl9AOcDKR
ap0XGHCfGqsvebVq2UPBpSRn+nFGoZK7/lfGawLW5YkG1JExl88Pn6cUq+zfafhFA76l6emL95DM
WDz573KU09Gz8F8xGcd4qBjgkiGKBmXUgDxP2KrNxOgiszH66YxLxj/Ic9LyTqbmFNS5dlwLGZ70
i8FjsIDUhuUbJO2XiNPxaw1YRJuBV8uh14Xv0Gb4pwoLHi8wm6BsuvOvAMnb90l9ziRR48uSbZpc
Aciwvk8rk6iyEx465vh4QyZE3wYpBohrLMdTNDO8oxOebR2fMLUQiWMUMC8ZhZ8th+dJIQM+8fz6
ZaLL7Xs3ShOWSNr79V24J88TM5TCwqLbVHyvgArgpuC3J/1MqM2tq8HcWRyxsiUsM7RAmHo42UQv
HsWuj61AVt1Rd4kR1BxmlAAYPoD5vmMzjYPh82CBZgIyGW1oa8TjdXOO12ylEvdeXMr82LNbuWtv
OwcEpeXWobzVDgQLkiAZ5KOHhB6ZNoaxRwof6qgBeMrVKfqJIKdYwe9LYW5c+WTcROFILuOoZrEi
DYcQ4BPSDxZMahgbwjsCxJIc73rpCsgEqlJan4ULoAkatdGBsbAzicUlKcS8pHj7qQqF7UKwEaaa
Y2MO22GmAuPvWZHDQ3RzCIMKVHUcm+tGzjZZi3XBPgxPeD66/RHTxwvyDlYLqB3d0JIoTV4jCNFu
ilhSA1vX8Z3I/mNEnmCOnbTaoXi2/ZwuKmYb17NwXUnV/a3QlhnxM/fyMixF49PEBmd8G+r7PuSe
zAfY1KyqoJtZRhyKWkRJ6aMlAczlypQ4L/8iDuNQFe7WkeeT1k5YeSWbjKAwvUIdQ4yP4eAyQXHr
Kjpnoqw4R9ti1x3/n2y8ViMji5fET7/inNN6q3dfrURAXWKDGMM2sQHV5RC1xMqB15FO5UgXIjhs
UtutR1jT0kPeirvLAV8Fs3dkMsp/qrsGVi2fvBhwoVBNzpyJ4GgJ01+pv+xIaD9mvcYECo7vEmOE
fOCjSUYgwHrzsj91iFZdWFXTgEkcXc6u1vzGY0ZijQ6FtpDxCyNzYj+Eb9v2ywCNtGOfxk8km0hv
E9aYUG7s7UfPmXEaSoybwBtuVUv+kUmpBuabx6zjA8zxKbFacAk5YAsotcQk/aBHq519mn7pc/T9
xb1+fntOsHYPXX2CAiFMMMzplHJMVjD3+Y70F96YcmgXCoA6xyNvrA6uDrSa4lcggPrah6iVr5Gc
aIqhi8ZRIVX7K16nCq6X2xw2YCXMndmXBOifJarz/yC1IwuBuVYPhMRwBX5hfqNNDNXzhPCs+6X+
+Cj1sqEnvmai7B1q2pXZ0AEOrmS5Jw3kxWXhvJKpNoInwYlpVCL1SsxT5xtY1VlVHezNsjyWbck4
i596N0/BstFLe79doVk30kiqaK6aZ+6oz78Nq3bXi0yPpdH/Bnjo0IK4bGq5Kg9Gud91ACcrvIFw
vz1xaT6B9OvHxmQY0ASJVAvCX4iIiMWprnW5BiK14zYW+ZIFDl7bM99E2DXxNRFzkwqlb/3PJWj9
EosN33nCjkY4jUS26sRngTV/7f02FLpoCdfQStpksZLZwDojLTHeLSpNjL9U3DhbP1OPMJ4oyxfa
+N67qX0wgmDhsA5/xjS1olr21X3pLDYqLjckcrPqJABQeTwxPCbZaf2r5BOQa51H3lNAFOAU+6pX
6U5JkEMMZmOQakSjW8CC3HcHPD5xvW7IZR6TUho58p7rCtwiOZnQHUUK0aG3R705y4D/U0bmSSQG
5v0+QnHNV0m71lkM9sAi5iDlQKTfyS9zC1LS7/rxxSuj3QtIofyk1icS50Zkyri0AipfkjUJKRZ1
9P6N1mzrkpGR4yY0QUDa1k5Ec02RxX0/YxpFHNug5XgHCUhuwDnYK+QBdq56RI01PHu1UOQw1EHJ
Z/8CuntrvsPwoPaMN/3duOy1hbA8kPApOr0aYRIDQ151UU3SrKHm+pZnW3ABQPMjVcmN8fnH99gk
+mrf2KtrdIV5BQVnuRoijQTcAOeH2OTSxHyTDLDM0JYyB+mXG0l3OWKKZ+xxX9nkjdNDb3jJQPAi
R2t/ny4IO2fjfETTZvACSZ29VDrcKYVhQVEs9Oh8214Zrl9nGjJ3xorJQHfFVjSZOYdPVZLGAcu2
cxw/3HenKmj5FWeGBihB38v2LVzwejSwiYyseMhs9aAi4DFgYBZfoJ9sfwuamP/Do9H0OpkKBUNa
l/Zj7W6H7S6NO2vZPvriNiXyxLl6Ps+XmfcAkISjoU2gRbwcqaJfheAj3jiDtYmpFg3pCkGRRqIt
gXNtlep7vMwGqHzOHGMwF3t1K4yDmrtIPCpYEdLmbMV2VZI/qEc6P61whNvv8VF8b8slFd+mXUXi
X8heNhWYSvSNn6hkPVLHN5imBEpPQeO46rKpXv7QYUT4c3i6MppHTBxTeggvhahHPAevWwZj9JTY
CIGtNMU9g9y9NBG5EZwPWyftpAb1Hl6303ToKo+96CcelphH+n6Cfxv8JSW/rSLIGESeu2YR0csH
5cbAtdbU6Cq3fWDBZXqGN1tS3EGC1Re8hvSV0GPrdMFdrJtXumD21r5yUMU/r/MkA4vGLo6Ae7HA
RkxOoGBYsxKf2+oLNNquDx/CpOJksmXYBE5UAy2RADTzctX2Lq/Kb+azIPIg8jzRtEKWJ72vTZOk
toEATNfVvIceuAalZzivo/VP/26WOhjHMR55odLdkLGJgnuobsQvP7YIGLsFZYFsfAiCMx05Jy1y
Mst0frek2ZmLDQtjtJLp2MFHcZmBeGa1kWIgo8GPxCuc+0asAykkBY0DylXREbOfGMRg6XE77zwn
m9ifYFipjDZwC0yDV+cSlhymD1H+4yoqGcvQnvSXkQniXatMwU4DELlyFqNMJs16NAESzNN1yQ65
CuqZ+aOtR6aJDlO76mQXkXw8z5E+3TiNH2xSSms8uDs/mNPhllAA3vT8RnhdbUDg1yv6eNUXlfld
dVVfplfXWj+ujCbP/PywIzlIRMD/VMOPn4OGcbsh7yiPnAhbC2zmWSjISHO//OvCL4GWILfRNdiB
grJWhiYxM2iMA+C9vt88aKxgblp8K1vCNpjola1AN+2gwJaVVCpsftKBJwnq7L+x5dt8fYr9fRDG
7Sseqj1+/ahb/k/FhC8+lOr22qL8hF2m8Nu7fNWNBp5Dle3H3IX3VYf3z7KJ6HSkdjx57arvpU/i
qqs9VYqRQ/XZE+Pg2dRG6bRgdhfQv4narwJGLL1nFc0roi5OgK4wfHMNu6Ie2PZhByiZEqieVLb/
yDqlrcCbL7EwzrJQxqEzw6KqhYqsH09sLgahjLGSNBqraxEEYc62hxo8SJZSGTUlZlG7tQVqvZjK
7o0MWR9jPgnD9a7TNX6q5nI2Xovdqqnmvik8Cnb9MUHjD+o1NGwLFwzWidih9v4uRaSFV7FTTIYO
AAWcBoa/iA/CUASC0VNJOvuWG19pANjDO76zLDBbsYazWfNTNLvc2YAH5c8IZDanA3YwrY+t6XLu
r4bE4hU1d8NClDenfPU49VApA45MSQrHSO74xrgRlR7W2vB9sgjgFBFPRvlbCrp3nlVV/k7jIVPh
cdPHC06Km6z9KZT7Z34ODtfQmkrZHu5LzrDr7wm/HlJHS8agfCuHQI9FAt71U66n2UFpIDdb8pAa
64HO3KOaGHU5beTv82UxizNFJQW5GkgwbjSDtP6eSRkK442I+PK0JGemCy1C4FP25lMhNrLZnYo2
8Q0y0s8/Z1HhQ+qs00QQxgkgsW3fG3Boq9WqZdaXZN4C4q+7kSAvEsTu2HZh9qFCxe5MgonFiIDH
s5IoPl8fFKk/7vKJesejSyBSi2Knu0geIct9pX6D6z7SRGS2zhxxYpYOb/0V2XgXInq2h5OtUO3W
W0XrGjBAZgSjrR8Fd1AM+aMdeJHxKRATmVcc6Yz6NmFPBSOCVD8Q9hfN0BmCU8u53e6kSWqm6wpl
au4MheBJHaTNZpywPEHLB693PZJkYg/I/YcqvCnhHhSk0Ym4OgBFjaz69ZbHuaogRdwg0Mafgd9C
CyfurNYW9mnLBnijkUotyCMElP6LCYWnsY3fMdHq4djQ6z0DbGD+n+0GacEBeGc+2Ovf7w1Fx6rp
O6Axca1N3V97YWfU6Nj8Mae0lT0iX+rPBrhM/p8NcRoffE7/lC0Q/kJ7HpTuqjWfzTS1ES8U6brA
LkV1GR+hHPb9Ow1NmuS/oeAYoFgFZGMQft1zQhs/YDQys5ftvpBJWdOK5t70NEr1kIRBIsyVto74
UhDABS7niNy8W4dq0+90AzMYtovMkSyrA7+Pk7Etf6S22uoP5MaukCOAZWAAU5iypIgRqwJDEXn4
/gb8yZxS4tBRJOBmeymKPyRN9CjykACkx8Z1Y9V/UdP3ZbwF+wDdq+bk/5RQ0Tc9QyU/H8ysGttA
kdg3yUf2S/MAr2E7x/Kiq39cLEi00BAH2EUjknI0tBeg9LaufIHv5FWto/o9L4+aTzXBJgLAH9z1
2wX8mhjncBXu0cpr64mot+NhuByv53C/V0r9dxMTlANuZibQTt8RzU18TfZCGe8f0w21ebZ5/44C
KBiPlgRMj8GymPbYplUN+1ihDITi3sug/jiRXyoB3K0pcX6f3Nbj4dKLwniRYAyfZzldXbjfa8OV
4QMi74/SIKYXwSoQupNyOOmOHW8gMTzTWuhpXh3OPvrEEeBUaYAcuRx8+1+sHb3qsEtouKeK1gXO
GCpeDLa5ibbc7bh7K8juo7HrCr9V1m5JxOIUh3AhN0hIxjSawVRJ/LOciP3cNDuc4kST64j5Qiao
1Dc5WPE3c3B8XE03Q2mHttPPin+IpkLEyjmxlCEEOe/yOIBvWbA4kQUguqEFLD0lFTmDKenIEp11
rQ7Nl4Iq1060jn+3Alb5nxzk6jnwYvwWEc4OTLnly29L/TqQjzqQhzlxvThzK8k2PStEoitUFend
dEqxNiDr0MY74t0Hkq3L4jC/pJiREj4wugSXhoTKLtwtkRP28d68B9rczudcJHtkN2EtNZJQ6V8i
ZZROnfM8Dcg6HbRnayl6rvHAh/ILOZspCv8Lpwe5Gv/UsnSz0ENPVMlA7yhBfzOLGy4pL8mMaGEB
Vp90goo+GL7INJAiSgLiy//VsquI5n6Vgn5DS3Xu6LNtHZWdnGWRquE0LpFPS39bEBPJ5XuLVhDT
crONBBFc9+QMsJcZJ17IZSjWRyzV5M9BfOWeU5fw/JDJl/FvFf3vm6Mt4a9XYgP0QH4/KwO24712
76caXcDl3uPWIHp1nKx0UfK3zr9tPxhXrPii+Y2XdQ4kDg/MQiNQWyyHBhFjrDxAWlVSowquebbo
3CceLA4Uu26eMYQT6F2Qmrs1S25icFpa59MVQtMEOFZWCb0QvR/rh4u2m2cYoeejE5t2BX4Povfo
OY4aOBwqPX/TEJzyeT4Q8uPPwvsFNXdTc9qQkhUIdsp0Byb5JsXAFeFm0TCrjrlE8gfFR9ktJG/+
aRbR1Ugeam2qX9cNfXiJxMPMnXIVPREA8e33oYFESbtZNMOWwkwfAFCDcrJ+xN3eOl/pUBYjyQv6
2yKzlvP0o0qSl9pqcXxGLR5dINqeyBoUMVLhKiZ82E0UDwoKZNWo5yU+IH+uzXrbB0pvjC2yiUwF
Ct7ZP2OcGNEMUlVlSfIlMJzLefsQkScldT22e/biRAHe5EmLqFOIZc/pPk9BP7YhMILEMIxYkEgP
8Y7xJ0Sj0MI+DWC/PvnFZz3hrWuMnD/Bnm1baGyv6d3LtWrqP3rrpt4rvDVHkg/XwlEmtpNV+KUT
bFklcImDoOj1ig+s3DfNvTS0zXjU5hdKVaqd+zM0DR68zTP2G1PtxKR/YPLhfpiYxW55IV4K9vyB
wcIXZsB4HVK94WrzsMOAdauVcN/pSLaGmHdz4Sr1MgxnQ/ubnzlSXVlQ7jXNqKI+oqAdMJBsDGEv
Vw0Sroxo4X+N8VGA+pePm0B+7MrCz4PHAdZcWPezTBZ9uYfwjl4cfLC2KktQElLN8uuIBlAjNTPs
+RxMqkqfMvpaYJdsSEYQ/AC1hmMJEt2P0VJp1gYbPY+Rd7cZDrEVCFL8QApNAxYQkZjtaQ8Zmz5M
/fd8E4bf4Y7dDa6Yc3nB7c0cadqasL93j7OJoQObemlaSsikcZR4/QZUAVgg6Tszvv84uI/bxJ2Y
ECeT88xscew5jVM/n7Of+5GD6s1u8+E0yiXxKwOGHwrJyIr++AuV1cmim36js8dALzh6w42XErbs
AwDlsZGsAUB/Jic8+yn7yRZdcv9AEnwcaFL4Zmqa+3+hSPrmaljFf61SG7z0GhlVnLY8y+ycAykB
TzzuAbvz/k/yOTdVZ2IUzYAB8+Hq/phLSjKi+fdDqJPsh+SHkJeRaF/QuplqNjn4GLKqLQ0NJY+6
TcamTn7+2df9IRvHeUJzi9Lep2yEYIL3m63Qp6t7k0gjRkpGp8NpmZbKervJzh4k490xDdkTOhz1
oe8wUyffl0W0mYy5yOtdozDYC4qeB17Cz6DAQUvTP4sBS51cIsB4Uz++er+VdFe9xR6QyGzl1GpF
YGOCt2BvgpVaYUTlJ8VNULmjK6+cBTiJoAuot7oSoaLSU//lD59q3Fvl9xPNb3sUtCKaDDND7ypF
82+uI/vwq0ZZHmOlEkeATV36/nqESCEOG+RiW3t5h8KwKZ/HTevm8epoFYegflNgyKeHzI8jUhSk
5dhRvm6ISp8TZd6/afr8mFThbsQeQu1Q1jq6wV3hLEbwq9TkJUbd1RmEqxIbKBP2gDhpIGXPg47J
QqG2znzS3ArB5feSNCAJ38r8SO/PelejWC+C2G04GSoMgx8aAAfX+WX05Kci2Urira+8KjIFKtjK
TLSOL2P29tFmXxetxZHUFpiPDCBc3QTcfYcfkOMutYoxe47uOaet2VqYIG0qQGCCXZNyL+3lOvT6
CWN4uogCWXv50yYVedCNFVYFqdjkISbWEpgyCQS34o+EjnOdDRPs4DW+Bi6+k4/Rnci1kSHoHOfL
UTleT0cDz1hQfnQkIYy9LoUZksz2zHV3jgQE2P7CT5GodE5eKu7mdYDBWR3GhygHFyo2o9Pl7gHH
e+kGlodsLEEZKFvHI1ZVMWqgAgYoBFbi0l6LDS6rwUuCn4Udu+Y8NujVFaZJZeL/A6+5F5OsQiSf
9W6L8zkaOsr5Xiay1Roj3SdebiAI9DMO9hhziSmtFmK3JrB0ItTfUFYGZRukn2HzsmRCheFz78cw
cFU9Yj6fHT/P3fg9M59rKMwmG4n53+3dWw7PXCAPH9pW+wNhaaPFfbUKeNToWqZ1F/nIzT0STRlI
1LxkW81vjjCIwBeCCiG9c+ziaHijjzv2IQgJezJTD+GcqR7j/3OfWQL9Joho91WtSrLo9E4JIyLy
fHtX5Kn7/JG1rQk/FduUnQQA9Ppy+dio1aDoXPxPYQ3RfgGNljT/lcQNN133Wc7Hcf5NDZWJOe8z
4C07nfM+IteerWvCxDVAVaCcyvEe4zSBo2eK13epdSH3FZSkHA3JRqVFxVp8L9FgllQL7lF61+jP
TwzEnzEIvk0EtmS8EPhbCZeCz/ZBI12cqSrEyC8Eq8ziVYWy++6yR72MBI5g/s+ZgIvF4AdH6P0X
SBUtaxODvnlUbKEKoKpmj3ilXaSRNdtjJNbQcN9ukDwXH5YY9Lr/m6B9Zs0h9AvpUpBM1WCqDeeu
x3voZENbHLZDa8L7IKS3jew+VRri/GyiyNGFXPez9A23Qm3KQKCuWPzdxERzgYA2g8uX9ZY1Eiz4
RPC35/mnzfKORx8g9ZaMZjrvu7huyULiJMhQAAPbCEvp7ZPeC6W4YgkNrQ8bmoanhtsQNhvguLQ6
bNBhkzeBA+ivu/3gAw1lPi/Qv1ael+coxx+YuUT49c1HTC5spYiHmf7VJo7Nvlqpw+2RIletai+e
Y5JF5rYdjtpW/x+qVQLiOzTO4Far6P/08vUtBEyUfR1C+0SmP1c5r5NB/ycrfhJLV8wOVF79xac9
pr7G7D3xzkT4fFjssuVRYKhJG18IOs+WIIcPOa+yaAo8Ro8ZGUmm5lf1lAmMy4p+YfRfmgBgDRgy
74sVLhOdRE+3wFTW8u7J5JB5f6t6KQ0NT5g1v2Te95NvtoWT6NaK/tHSAOMOTzuur+2fLDGneOjC
zgWOxQ1kYlSun5MIdEy+BrMRbqXt6dk4+oRlNiGSC3slYxR6fMWG+1BOz3OiCrc043RLwQb36Ioz
CHhQMeMV3Jq/vh/qMPbky3Jajks7/Wvh7OOSvEaIotR3RWzAF8IvFD9SRGsCdLCxHLoHVL1PuSZ4
ybuTxLmnaV0gdaO/VdoS2KqXEtTYHjW7LyApAMT4i3KMtZPoFdfFxtd0MaMjEYRjnnoDesKwLtIg
3Gl75b9dTU9M6dr6q32hJIxzUOuHnCM8aEArH8IemaK1OzeZg4ncqKMBSJSKb/Qcg1JrOvrMNMcO
pMiGDrVR0x3RzkziYZi0Q7Maz3v7tB401o9KDpzikmnOIYEdf350Ku+4cgZ33lwmlEf37wkvKam+
JRS4yjAfNtm/KTzm5R4pr4RttpoDY6NUF27nUSG5Zx0nt+ibCOAPv0VL4PYVf+CuRkkrRtuDjRCP
yOfu6pWcd0U5Ix5FcTc2wpSPA807R1IuRmxXSDTQKrVCrLo5idsc8u/nMOjY7JvdIfyYh1mn47u4
TXNylqfXPnlJWlBR4/wgxcbFnf5WZHvpzKLhWOlZnqbYnGNDjc1FlXZoq7N/MfMFqg6CAOBChe4m
yaa3OiRl/LpaTPB3ZuEO4YydkM2z0H/2HrA7Qvfqj7JyCKKwabHZ4na+HSRw0QqNKz8GsKw/56Zw
IfLq9FZXkbf4EDZTm1TCBPR/YeereIvdoD7pgF+UNwuat+GntSFQkIlE9PzndOb66iHblhwLJ9ri
+ELnEmewFEJWRZXpq0+COjEJqoiUOqu7hCFWMon66MOeZRNDBD/mSBu7fawNXusJ1PR+4GFRZmjS
JIeRcCCFM9nhogxSNdNcTJsAleI97Zo5muWkfHp43orxgwjnDdhz1rHH1p5GRxATC69CN2tcEZfY
tqh0G0MlbJPP3S4s33llo3K6ZgG/tPselgh5jBnXRHvDP5D5dFeGDgy7GrRxcDNVMQDPeRCMRR+O
CXxTUXdneFicoyUuIlPKQUy5offY4mkPZ2a1sz6z9GAqJoryvHz37HoBdYniP0moVlMUiKBY/JKc
sTCU72xdh9IHQa0JGwY4NgxRam4+DzUKr8XZh9CaVgl9euSDemOuRpRcBht8q8uLQt9nNNwRNwBm
Gllsos0tBX+hJ4A5OXBkcbNNVVJiOI8C7EVpVSX2OtDyHoDsM+BzTwCGen4OwuUBq3VRdAY9TcyF
BJ+3hKEwrJp1M4uMMcaem0DZpZ9SfItHgY1WjWELkrMNj5JBXLOy6IdVJKElkjV80QaTkx4KKEA6
DdufOxpe15vJZx0Nhj4BVwwvhV6b0mRRr2RrVu9PxGytLwBdTkK87omR8YRfIcDILUu6Xn5HK3fW
ecvJFqZXNNtOoaSHf7xaftwvPdnIMiehzoAFpgIetkudDjgkup2zHI5Xi0n4SDr7b6zo8hMXp9Dm
Y6mgRJHrveh4l7LABM1OKei0fwiOZWI3No/ULNFPXuUEPbILP0YSonWR1nkvMBb2+OzaOsxGun4w
n+B2YsKSyM6tPfAnl/BMuppOgv8MWVmme4K389YdI+hrzVRw3gCxolIq+h0Z7giKwqNz/dmNe0/f
4MBdQSrxX8y6f9okvejfVyei9wyC4PdBOv26bCvj3mqt8jspmhERCgAh1B/vqCSfKA6HxZt/gn5/
DQA3UrwLZMHyYcopPXBkKfogqD+IFry1paM5kTZyAI6/ERW4dEJ/1CtDLYiD07LWMYYi/iTtLHFy
6uwp9fQ244RZpWBqgQgoU1EVUfcPe70o30AjqM3UALg6Jduu5dol92Lwm5mBtGLonak2ANSsMJTc
HmoQazHSjIA6OFY9Yw8IkRGZAVfhtCSbfQYfaXfPCDggW2BI1yBEFlmmDN19+LZoFb1hCnr+h37k
78jvM2Bc0m3PxvyuRoijoC6+1PzXykpwGAwgUoOrD3/hUYOqMWfLhWdIeNTZwEKaxH4YSfC5lXJl
pUJVOc7cWy3Ss07eL74+UGX6I8JfU92B9fWAoKx1r39OK1jjVVc9MupoT3w1331sGcpI0WiwSUdm
SOv0kdPwTkZBOJXbnxPx59R31RwWT31Hh7K8zZBIbckF+zjqGpYj4z78w771GthcH+SZlfYo7gp8
Ri85zrxylpe9z2+AuEceMmZxVqb1dzjtUrdbWsMT8vYWonbBBi8HjI9aWUwG8tW9q7EmuvosNYv+
T1JA+MsZiVrfhXBFqQw77zYZgZcQPMxJvG7ncFPbPcbaIG8zzK/tCpm38By83u7igudanwg1E0AZ
nOfja+i05cSxcvjpXer6S69gTfSArIUUmWLV4No0a37AEBeDTZ8sgj6cwq/N33BFWksz8VLMJnn/
3BQIav1Dp2fg2KEEDvno9up3PnlduZGVVkLD67/RiJrv8x+1++RKMI6IwpZYeHapPKF9p9PCIlO4
TGLruIotZtkiVFTHwokx08Uxttj4076CKRS6hUH/9+e9+92A+ofMzBP2sz4p/gKigBVELmfR80ht
oRGFaM9aXDJantHnPSCYg+ne9x/ZhR25vjrLUhbhYR42rgPqocmDRGV2B21Z27Stx7hB+EXeplgO
GKHmYI6vDzG7VWBLQgNplknWF1xwjpvz1h3py4WoT3+KstR6qV7wkxMaJRn0TataIA5bo/clldgB
aldSRaxkfiTe5mhPaWCHEpzEWEW9AMI8pUD2ZLo/NP0LUr7oYzh8EJEswWGlyE1SUrLCkwZeUyCo
Lf9WwjqYpUC/OkrCzNNAR0UN3WtlbLaG5tGndsETX+C2GxP5JwKOEVUv5PY6VaUeE41VnjaHVUb0
8hm2rBoXQmFNCJ68YuIoeYtKBmnW2Bo+QipL/foCsh2OZ/8T9OOAjyPxdg3oFQYvTMU8fdR0aPPg
kcDw3dK2/S/UjvbKROc16Kxo3s0cKHU2+KHyzdoWnfQZYHnZyZ+y5WiLJuVtavr9E9n2c1Rzm2Ia
udmerLqxPzghUd07V8lxk3wnnXcBOXVcPr9EUJP6mzFRlpahCxi4pBprCtfscsyFvWZVEy0tWLqX
VLtLnXdESKYLf/MIw0l63Avrc8Jgrnyq9uYnnXpvVisgLjeDp23Erup8sCuH+St2OW9TkKx/I8h8
cLvKZK6N6f7X9TGLUmdJ3tMbqiGbNwM7nhiNVJfBgAmb5po2vG4VlF5NawK5DYXXtUUXx2d7468Z
PSWTDURxMLUjD5mKiipN0oNxENNxjutV6OWWmC3ksKIrMMfvJpCSkASt42GMha9I9QmqWkPJKx5V
NxNViJrV/n0VaeWuXQBI6+V5Bs8Moq144ESO7AfinTxcfrWLwNNua9WJXbWRhSYNcsPGcQFXxBuH
ABiwtpSlRNTP1Ft0PFxenlyanFkkNMlLR8YfmoBfneL1T/VxrxkAMQxJGFcUzYZVQXS7EHFrWqye
NjgSQ1yvLyZgEGCWXcmi3K2Wf2NBXxV38DRX18tkzscraui0Buw10MGkqm3SqyVzumieBGNkVRaJ
QdLk7au1eR77PwBr74FKMedbLi0h0vdqBmBbYhGY0T/Nfu4nCpp3RxpYBwsYrwVFTTgV8rlFCj2f
XEk1lKMofjyKLMtMdyJRs/gFeahDjfT0NUGUAg8sAcO6HemNynSVuwpZzqkyU2Gn42cb6++Mw/G/
gyB2zjV3v9YfYUNItoS1IQ6Rl4aLFR+4w3Ndfc4OZCOMZjiIIwsugpg42HcJTsIjSTUC/2M5iHij
N/++Lgm3bDaElSSMzCei7tUaGLoY2Yidzw+/C84nhxlEFNGhNcVMYqLQ/xsU9nUvIuOKuGCEjk2c
CAAoRUYYMXug6DO3ujlYvSXq1SaemE+Tsi1nQkUP2U6m3JbcXXFkRUYT+JmYj+ao4Qw8VzudA3Dk
Kh6sYwp+OYa2xMMsYpNsLT9HzeeNbPZKKXMWQMHsYdbpj4GnefKZJnluGwauJZ9e6AvWUoRTFdNQ
qYeUu+z5pfIZnUrauNIvcRfjaa5fE9RMun90sB2BU6Tt0n87KxHcn9UAhoyeSu0tfQFAFQm4hwfw
M2hUE7t2PWidmGk8+TVQDFDMJC1kIhm94ej4ZvE/a9RD8KhQ5TNmU99l3SLKsQXf0gI9ZD6hFGLn
oNnWlo5TRVN9wPFcp+YbCjjLH0EHC/8I+marGrzFiqUIQ7NDlyAKxrDvjaybAXPcPob/7GnkD0Q6
844y+fgmWjIGH+HoqBlBtAUkCv7gRE9VrulGt2prP2K9eCVRQRzB8+xPeJInb1FGroxgWDe+zol4
K70seBavFhmHR95y10EDMa75BRo8b4JdXbH/6CMzIQen9lZwsPV21lc0LPN2UoS0bLuuaHVG3JX2
Mlb2WX6b5zn3TzWFPSx+Km6oNN6F80s1uN1aeMT9Cdry1c5jGKf6NIuUneqfFlsmf1CR3ul98ixE
NVS7gZgQ8RjG1xQHtB3l59dHozaJSshar6cRLMGd94j796wOFEbAC81tB3dbzhjfjJ6EGuoCQDJE
k8awBb8cFzq3Dib1VHqt4l3dmYKjMcPexnivaymKAhjKNi0BtXxbYD0yo8nK6mKOE3MX2nEsDMrz
kMzWfqwmMPWU38xGKY+MhEiIDAErP+FFtg5YFd7C2DD3dWa/2603zmGNnR7pN+Jk3ER0BSKyeK/R
PKaaanVjQD6MmcDg4T6IlAXQ9RW1H3+B9G3Obk0ZH+k7zfTFSv3/sFxDIzfWo3Ti/gosD5KdkTV1
xZ/mDn24/ykhqGU/Jm8FqgdbB5YEj2Qur2Os+FR33jilKi6/sKlRWgjNgBCR8rtpUCJYh6jEBgXz
QjGisxdQ6mPSNc3Xfk6YQHEoB1bApRoglj7FIKHYnK2D0Kro9+Zr4uD6DIhEGwrwavrJVB4/Bu9Z
5GYxAmNpFFkolkE1JF7vHImPvZIxtOTYltINxH2dk3C8Xgr2hTyuHTkmbDrLvjWAFoSRphJJlCyy
wVduX0dTEySlkGZ9Ns07gyO7dFZZyr3a9+N21Q4rvWp6A/k7+IURS0MIKLym+a4QaZXSgq0cZcNR
NwVw7LjItK1gvZhbqIxmyNDMSxNoz6JnRetNq/SJ2hoVoIAUFjhV7A1mm3DsXgn0CeWgKUTveMbO
Mr644j89pCvIqg4WIZva+Z250gIwSYTTgZh25dLhcaEqsW6bJz+Ktmhr5K+J6ngt+FEqFTwhj7eR
H9Mr4aB0XgFcKvg+lHUzlIloXr6f0QYHsfUNGLt6fxN54JztgKNj1UgFUQzWg0Nb2jTYLRQ9l97X
PuMymdEsw6K+RcB3JXzRaCUfSnzNzFhhR7jNjv7dS0BqeLxx88vQv4KdRwEwWCSZqwBJIutR5SbR
hmqXzFcQCAQVAckAL4gj10a5gATST2QZ1GN+FyoC73wKyBAJyEHcIN2FmbVbQkdv1sLYTEqU4vw9
yZQFth8QahYZkuWnL3AcyJpQtu1a8WFPo8/4jd1p8cKgw3H3sLcRTb5EhungeQh/m049UmnxFDza
V1qV1F8DhH/TeRrgPpgLoSTme0LnvKAYzlf2maPY7mwKOE14tP8YeEXYlpMNzHHMwT4CKHPNzieH
nFI3OdSU4et8BPClY/MnWJgwNBvNm7Ropb07E8752RcpZvqfm7bO2Rvgg7pTg4PoNjFiH8fCkQ/a
WzwBbaD+l4u4czbGrk0yk6Jc8yrJ6R6HJ9TzAMItka0IqIBCuifny+Zb/lnt1ASuWpI0ZC7FqKt9
HWemH2KX+nc3ebsNIhnky4Y5oMwWCwFE1vD7tDKNu3ebJMcxWsnaIilPLb89W5Q8m+H0A8BUWVB3
kwfvE2IZCxIkXBn9rntR778hEwML0M69PIKRnFs0hsy4maPFvDCbSy2NZYMio6jkdUwrNFBcvggn
Zvh3yU9BxPOjzK4W5rzwKTF1tKzkBYi1rjjbjo3sRVuo3SIUh1F27fWz0FAuSJ4QGjI0kpcQgULu
algCB/kA6QKEXD7nR97EXK2nIvzyAOfasx8Q7cjixwK5S3jSfLy2pSdOaQ0nR0KEfHmPNajvKd/a
Fapq5vjOKQ5D+ERK1dyR8enbj92RIqYKA4PdeTekdNiJ03fY8bw1ce0UYbStoq+7k9pF9oxrGuLy
t8uwOs8R25P+I3KYC0qSsPmllLGtCTJXkx9NxCCZFwvLPzPtn+kxRLRN1qCSltrUTw0kUITZ24xo
fhcpgNoJlCzatISyBSh+TqektE9IytpFcFNg8rF0eSakodgtsovGa+sFKJ5pm+E6289YTMeH5Zt1
Rv/kW/n10qr8De4VXDkt67uCJvHsAaSgrwK8QGu8g49okSPtniAm3TnenpP+ntcOHsnOEsiq+Zru
8F0SBNBo/p7rfNfHv0qSA4AIcvOmMW9gv1gSmSNAXEmoDRIWgT8B45UBJLgeZtr/83MDvfJbUPTK
Tzt7FqpyrKy7w0NkuRheg/ErzeohDPDTBDMO8UDHB6ksNwnUs9gaPTZJ4UsNVD3KdBXmKOF5XlJK
gzQ0Hmn05GFpA+8WaNa2ZzyP11tcpGRoXdbR6Bb9WZH6LIOfCWG6062vfZsiS3If+g/gnrj29OA5
9ZABRpQzUGFqx6Ecy5Egm0+DcueYLAlVAsRAmh0w3dSAipPlMbCToc1bHE0/cwoxJFYuWkkDHy5f
CbEsUxFwQf3cl/wNj4eJ24vh8Cr+uq6JqGzkj0HcdNHDyj88jHzuXbo9nJjr4MgNkm9s+6gDoK5u
px8cwizZPVPfrr5XrktUme34I9UtI46vwE9hHuj++6jcVHnOAf9jnoTPbUZuARyKEdnNCZRXlhQz
u7ERFOij6yKbfNRdUt1sygZQI5T8DuNxZVWGo/cbHBYK/fD8RIOVZAkrY0IadTwxsCUa0gmKKpNo
J1eIi0Ald9pIcjY4L2GgfPWAbMhhkSrukOrhqQ+/d2iBzh10Vm6pfsoZPIx5JSN5h+eMqxr63hFj
dv11eTxCZ+dDe3yRFDfQPZHMDmjj7V2tI/DboJEhWWwJ4Tx6zO8kAd+4//hsijDHLUSS+LMdaj/S
U5tqaamJv4DTaUvSDAlztWekEl38XgcFlsndKea/DYRfaUVF/Yjv+D1cjjPzKD0PGW2IcKqJWZji
WEFmMl/DKAw7
`pragma protect end_protected
