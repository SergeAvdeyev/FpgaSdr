-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Zqn0nzStCV5F6wGUT5cmjay5nerIs1UObqmK3GOYXwuPTfL6nqNBPsejhyUqQ5HEBCLh3cha3rvD
xdUz4C+0Q9nOA/yxxlhjWTC6e0rnRhKLyFVXheCucsyUxpoAIpoktSkRoOUwIhaKpldrQscyHoKt
RiV2olg7PMXnKQzQYfuzo9qFaRAst71N9RMUqlCwMBgYqGqrCRK89v2Ksf8iLTN6wOrNVfizp1m8
QEETJQAh6atC6ndS9uK5nZhALomtmz/YK4RDqi3YgBwP0p4tslUohUrlFFkKx3+M4+TVmNMZ7K/y
rMIFnLTxxGVTqm5X4Fl8KACX7KMsBwPOxckVmQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
uyE6NvnIqHNzvGnJvYxm5K8XRUNMi0EZmvlOJx56wI1z0LmwxDKEWswB+5FhTTqteSwNWqSDK8uL
DhoEUuDr37uE2jlAsavtHBQe6ovmPJtq0E48KzEXjzTggXEy6degti8k8uBLSUOgI+KrB4B8hnEt
pXryh4pNAhWXkZ2wOUvAyf1y4nOc7jYZxhfebvrwyy3TOdSppHtDdAQv9MZuV8VQy6wpe2sqH6GV
PDUQuo9Mcn4XNjcd61ZyABXhgugTBIR1XrZSEhFy6KFED3jmd563iZLlDnaH0j1ukl3JxCmqt7Nw
jePM/QVCsWwuT1hcLk1jZ2NTYUOQMKetRCxVS+P0BL/YWr1li6R32yYeeU1+RsydsNCC6uTrHYcg
1bo5mfgbTDbnJocuFBFv46di44vBlEoMaLf/6KQ/99v6Li8/iPtgWMo3jILr+Rm3LByMYsnn5tfH
X+O+FWSzuPEL0E6iXZOwtF5Opj+nEcuwcudtDQ4fCnd/KMjmd4zMzn+sfVrDmpUGWfkMUfprWD4y
TbMndMuLwp/cWpZl9xui1xxjPM1mzbYMxsBRy7mwkN+2o1y8JrzPFe6aG8cR/ugIXBjTiM6/C7v3
ANef2UNppCjLUGpnMrby6PqGCo6jqqpDhHi9uS/nhxfZ9/ULfbWE8b6gHRps4kDOPa6u5E98woea
WLKl10yI6/6WuT0VUaPFJV2Fr33bnvJi9t41/7aSItsGdyIsK+czwLVNKmYtOF9EfdGf2sFC54t/
mJVACNTi4x+bxVGX0tyLxcVCVUgOf9Ku5rGssasi6vb4+/G+8u03SRuzrg8pGcMHjWYCsfzhc1d8
4UCq7WsG5kUufNEGMDTzgQ8d9SNcHda/l/5peLNF7tkdg6UESsHjSQknreGFzl7F6WeDVPeAn9nc
WBqzHh4rVl2GhIP15aai/4SJfAmu7oOmKc7uIrzXejcvg3hhMu3FP5JUUpilYAuQU3IUqYYiFfGp
4Ne0ju/Xd/+qOx473xjFKgr9kk44WHRhdW5gqxc/Jc9EJuob/Hs4au6M9PBFOqJsmsfPcdVh8+sq
GHhorGW97zWMz9gKV2bD4grD3IcXX2Gnct4256UYR5aBrIb8JuIT8JE136gLfp3OBLRcxAhz/0XQ
bT++HmN7OqoqHEufDI47cMnJEkyaWwqauj4uBtHcVNpUmc8l/zVroO4j2I5rCemlGfE4tgcwKcyO
KVK5543zdErDzGF7d2jxQlcpk4oZROzwAEXq8rFgp6ug1jXc3Sv/QtPJNzIa1ncXSfBgHx/rATr8
Mnw1y9Dk+jEIcyEvBoXZogm4F8LhU4ofUMmZp2lTmeNEsQ+bUrZxeKRKXYBY4CqFBuCLGLjE/W4K
1Qkyk0allfoOFRpmRLEwvxUZzrOeLGpiiHVF8eTAwft5/9Zj1WaKFDgfzb7xSdsZePgsVTgaxVr5
VGn/XXfuBWz67UrWACy53DZ5hb4TUJ99kFA1WqbXWTOGelP7ZnhvzoooEMgnpFDPdtMwouCithUL
2utgVsen8O+1B6qI0DNA3GwATqHdFJBDJSslb/D8HWCRge6ScTJinvo9G1y9B9lPGb1ljlYpJhI/
6ujJCg3EArORDpz2Yn+zcsOCP6hsEkeBFk+1jXrxbPaQGg09P27DQ4ScQdLjC0K1abq/apYstQ8J
Qk35bcf1QP647rflL8AHwsOTid5R+EPLUwHRlrGdfcCSlXnlaJwNTmBEphxTqhhKlgE1KDjWz2+H
Fgi5CIWM+/9EpTIZmm3ImlOWXIPGMH6EU/FfgAA9jNsPFuqfRwz8KFoWSB5xk84lKS19ZavxuS50
kkbhcHtoeyYhtBWnbCIZIkEivRZF0MuDgWefYWXiljYLlbUyhcmapQQr96hsaAJ73iuip2y89w1O
yXZbI4DeZV6K9uJIRcb4GpdbD6Guwny2VDUV9ifgnxr2cUGpx78CSLnOLyEZXI8Bm1Df/UHgMsWu
ZcsY2O04SQt43gimUIbni3zUmXqRlJOx58xWo/bPsxrzHcJZoG85YKm2nxz1EjLSjqyO7DVmeDTV
AOIhRzE1pHMxldq7AUCtzQrIy/qMkwZ4N0bcJ/qGzvVMTzcEJor+XLHuZ1nSQJzjhy1gy/zTJ9L0
Zzl3dgisfLOUpPZoLFwwljS+U1qIf2g/cXyCvKM3zdFwvt8kQieeqwClKZnGSNYxXXentSZCEVuC
QIZ5skZ90ry6d5v5ghzYjTEA5CW2PFmBhQJmg/F3U5luAdtxuuiyMiLzRtsqvGH7HW97e9pTPaSz
VlAubZkghDysvNdVRL9akQAeKDwVdfgDcBagbcxozgRIy3cm/ERw5JkI0DgLd5FQgLsbKEB8Pw/r
PuU5wqZESIJ343SVaT6nbSsnCr+bcZbWhJpzHsySJ/XWa73wYd+I7hRhJCXrvOUviDl9d3RC6gE+
MFuim13vO7+AR4KhyzjANOWH7l69bmKjZgfQGDW0cn1UEICwSFVGMeo4gudOQIfmfzs9XjAhPYj+
lkpahizZAx+KVTgvCEKs9Sk8vhAqAVM4rkylz9Cselgzcry8OfG6kta9EfdhW286sRbxyfi8Q4QW
O85CuVFfv13GcZrnrtBVY87dMCJinefRl6sMM7swYGr+bGGnpjD7YMvwOG0Uwbg6k1EMA/bRWMgk
HS0WrxDblEpVveUSYm62z0cWHSYUcSD3srM8qabY63UPmVASjrN1nekgJcQFFmlYvXjl+V5o4+IP
gvtLgD9iwsgqWQgck0SyytuW2PygE7EzZeWihwyf544mHnToQOV5oT7H5dfkdWr5vkNHxu11rDcp
cMCKWh/gSOoZmRD1orIUT3CtYgveYIO6CAYnF1DcrekVimL8cWVd9nGSiNOWxO4KiLtKR4iJ/329
VA1bwj62XLe+ClB2YEWJUm2Z5Wu0cJuTiNWA9WfKQYho4+Hg9/m0QuTbG+6FNi1kwc4i1AWJ7dAh
f62P7ENc94n242f2CFpjAt1BcVdltDOcsDMzP7UVoC1fkB8POQkVemDqo+rhhO2doLv3yD2NLhyw
SV9eIBP1ls1XslJsMEAcK5zAmalSsbuKCi+UdpiDb1znAitNQ43oQdmOma0aAd2bGZ0OrWjXAsHb
3NTD5claaQPrYH30nlSMTdRykFjp5TIHsV+Slj5gergpZLQPFkLt206schVy5Z9uEB2yFqQQGmOF
lJsnJKn2RBOFFqmkj5+Jw4ztsjAzddWCj60bXLmYp9MmvRqbPZbO+WnY8Gm9yjR8tTFuwLX0y/d4
j4W5A9AdZ+dqM31hmnK0sZjnSG3da5bDlyuwA6cfLjo0eX0JlV+KcU5RDOiDSJbEV/nItgHt65mQ
KIqGiZaUKUUrdYewxs+fIDx6PofkpnwqBG693HCY+4zOZIw0Dhg4HnxagtlhqwKjOweW6M/Nn+W/
KyYUvCCJl0T6HKfPxiivBge1f0OZPzfQXartle0JcP4p6rtdmly8eLXnJtDbYmJADkEz5sLntCLA
mLAK85RLIA+1t5AnWmDA5oe9bw9w7IPCQMxORg/I+K5Y0rG/mtMsmbJDwYjERIsK6DQjWY6eFzmR
WQy33Z8CUuKEjWSykcEspCdBeyOqeW0XiBYXo3clnUwY5VdvERefmX669qtE6rDyIzeMp3nFVOf6
lSepSFMBQ16VKAlmtDv/ORlET3ZzYqxIL0pHnZ94joT/9CjjrVtyX6WXYqNaWzXt9LbltzogVfiw
rPUB/H3Y4hlRKfIU5DmmkvqvcCLVDtN6qUX5HGV3qRx6j9C9wfGdEW95EsvJWKCMMQ4lIOccZHHa
xS0FsQdDJcClJTs4bX5bMfd9BJNUYy8M0mfj0cgTIIXuWkPbKYSVxiEHEoYI+Hf4iF1gWAIY2NC3
CArn5p474v250abv8jrx9E4E8zTrFZvEFvMolAq5I0pvoPuQ12cAtZY3dGKXGlu4F8z/yiXQGg7A
WH7cLOzlwAL1mDhw+9OrWY8xmPWAoCBIIzwGsn3RXkJkV/WjpHLD5tpbzb81t3vrJOPDduflLG4Q
Bcm0U7TfIuivnzq41ttuy1CF2+11O2x8iQWPqYqM1Av2MOgSsbd7YshdXAJNtrGler/TDOpTKBIn
n8VQ5Gbu3lQmn4xbDBA5uUopl1tq/2HvC+XW6etIW4CamgxNf09h6Di1URyEDPZO8tDJK2M1r9X3
sbnmrXkArf0iEassM82LLIdoR9lvwaJw8h8Y3rwTWC7StnGIBrwzOULMijblT2KpRYNv+MC1jYgi
tgfGm9GxEtZhx2Wj6me9jEkDJ3RBShKOeXYTAKvXI00b6cjhg8ef/fe0spoda3DpK+zkZ3WDhfp+
Ad8eRm6WM+yDokTItjB3SCZjZiz/xBct83wUj1WlwsUzzS1cudXntAqVzINI0EzldyH0Tq+C4g1N
dcyfnWAYO95txS1d7+amITWycsnGLzc0C/3/uhCUB0N+zxGzaXwsHQiPkY0zXkVajAslbKGAf8wS
gEcLZ7Vg3/NA5J7utoWd7tDE1ZG84tbd4LAri4VYAu2zCfxSsk0U9j8GPjL6TZJZL/jjsZ2Q49U1
CLII34bM8u4mG1pmODQ/mDRGdm7/4tYshJG7mG2mYg80iE+R2VzOpsCTK+cdSzHTpsOuIsjnl6qE
WTOp+ySBketKdojA0qo/JTl4npeCdsHJGJX7ODAVAfB9/n0D7OQx2GvKSz2JpLIPvlCdnQroY7it
0r1CCaFeJd6abmGU00apnOJJSXSg8z0T3r+LW7VFm/WFqBuGtMgw9QvH22O+eFYntIpNeeHUPKs7
LFGXDFHoD31ENuvnrxpd21OK9e659fX8kIkJV7Ice2HhktstjMBtpyJI5nXaoPeIF1CU+aQB4shC
4gS9EhIatAfowQo1XyrAlM/Mnq93V1FYlIagb83HXHnnd8X0JZcRPZVj2QEn+/wAlJ39CExF1HwV
dif4hCiGOZNC2XP7fihM2r1bnhC/1vm0NWGXISuZz9PQjXig4/YNjqqg9kWoZb/v6xatHYyrEm0b
E1PZuox14mUociJLw1Wuz3KIXjj457aDxq6gKLjN6tOa9GTHlWvM1QMQ4RWku/K2gE3VMVY2HBE4
ApBQH3cd6yl8gKJphcMATT38dsOwPA6HmZgWfIRQk8TsiOr2dBvpaTRfxeK3r+RlPfuPRQdVQIcm
k2nJ/673eK60MNjvzMalL6+agnqNiBEe4cczqZJ3fEVXE+kMMiOpb85U4KfcHWiWL5SAmGJ416QE
P/0zY17cuolYFQDHMfhymyYkU5hLa1j5FurCVjDHKOEFQfKq6wLlyrAPjdbhQh4RisERjf8t7M3a
KC+OtAn8PzdW1GFStRhCx/xuYZHjADIuHEGMRvMKxnZ2PS3G4VLmV/N9OOpUoyhwKGzz4kKqIpM1
cVONhLkZRkWW5ZET1orJ6NKzHVTLfWHTlFEFkJriB807mne47Xw3htUpAk6EwoG0+z//BNtVOeVz
h+7YfVbyPWta8D4GqYbfXkP7pn2bXoNg+iVB3YPu4qWU78kUWxirXOesAJx4WduImAicS03JhHpG
shQiAbf6XgxGe37GRBLXCZ5MJ7C9dXrnYGOb/XX/RPerWirFvOkMHKiTwQuXUr3dcy0CqI/sZtX1
u++IEUMtZWljSAtIdrgU+eYO+3ssEZlpN8KZYdHoBaYclj14Dljfjy+/kP75oKqe3nYSL8+7coMm
fpebQrW3j766nowKB81jgPVWuH6LbFxxbXRbvPOjbULrW1A2LUO0ywjZK2YdNl8ojm8ujrn6BdSL
71klgB05Ssw6PGr69taedvDrBGiaDO0RniebY9pjGA9mtwd/L92+KBM5mlUAoLYbqPDQ/ThnVIHw
r7Y5Zfp0V3OqGtpEuRUikLJjUef6kAwU07DRhMgW/tVuwwKBGEmCLlmCzH/jXLVOeU8KWJ2rAeIt
4weRl0O8ORI/9puDJyVgjQnd2ao/JxwrhbnxSlF/HM9wdDdJOjP3EcG/LYxT9nsH0XJ4HL+FMW5W
Sitmwp6qAe4Q1UZ0FTnyiX8BUDCEP08zKBqHcg0O/W8Ibssl8k2fKhApdvVNFU/tKeMKplKYM0eD
oe4U3/xHoZe3LtFtmxNmwDnJ2uLxe1KYt/cHXRj2F1AgGQagV+TkP65agLN0jk3nR0oE8DVFs+bE
I9I6nEuZ80TwCDBITpc8yY6p6Xa6xPxO6vbJKmRTc5uTfi03q9DqPkLNLk6KxPZpAEdSqwfuHosm
uoXS6lIu7CZP+QCyjLOI0XQX0nx6qfBOoS1pC4eS5nEPxnn6yRUF0FGnYhvhHLjYhF4IpUK59kTN
s1t5FQrJ1jfeqCe7n9gvR13+1xrVYaRQ2yxv5ARVivl1xTP5LIzjI35jv8aeCsEvMxGuK1fwKOeF
r2HJomh9sC4oS1wZRyF/5G/Jt5drt38VzAXe5y07Xd2TYWYzOxzNivNpif6S+ScBtnT/3C5olWaZ
ho5LZfeGQSACUyUyd5YvHkL4sHsDsTrZzsNh1R5gCbk0T81AdFglweCY1jcQ6/IZI3zMILkgQsG0
APlrhVqAKQv+ERxblHTHUX5Rh4U+amUPhynsvdi4YJ1/R05PdqRGvC4EXzmyFopxGu33w+eQVDq+
jfCd98686aqrq9BthZesvkmfk7MJcrnytGIwWq8WjmrNKXyPH/EySzIVMvuoiz2OtxMFatXMXzNS
1ChoxDQLzuUi9vl8tpD93Gxhhyzb2lC8jE0L6dyvP2EQZa7O3BK2peNLEoFL2x5V7FQNK25Ly9Uv
JP3fWVQgdKZXY1Dot7WkYgMJ2ZguVNIzCfrUf6rhzodYK/ce0FNU85aly+hO7loKPi+DzzkiqJ68
p3KYk9YM8f5Z47CTHqcpff1+GPsjYjTGmzXZdG4B0S9GaxBfUGrZV6rsMyCkRrmmsGGpHLFJlkvE
PVzzhT8PudWaPP7PlJpa2ZVbLdFihZBXIHbZg8V9TqPFVAqf1YnkOcNN/s7HC8jkmdd2rv/PmIAa
K3hIVDqS1rjFkBf29BiMx3UBBdvHKUr8X4t+hd7HFZ1swUBNXgsyQUra9fIVNU3D751cBB5zp6sd
0xr0iSVoaC0sCHiBbi1CHsuq5x+Wz8XZsamtqtSgEl8nnr7LA3qncARj7j+SVAKb/naby5xz9DPt
AESsVNw6la5LhQp0l2OjnwdOh+9x1bxRHawRx442vFlsPQg3rL1Ol6JplCZHilLkhdyi5N9NXG1N
V5/G1DK905VgQQhf0FlcVdCAn7Ng/IE5tesu5N3p/aN6yL2I2B5DEZk3icJM05B1xtS5TuzUC+/R
61Kv6Nx5ORrh1tkJkfrxom6SnTQ0iZwFGry1ZNMYEPBwhOpvh2D/UhzITU1xGz1sRs7zfYVO5y7m
JqNwdDN14mNeLSfEkzkRKVhaCHCDcoPBoGehIZ7c4DZKAhatOGYC998xWQ5FVOlUcyB4vXgj/GJd
FgBzz++eWkdUKokEaXiK81aB2yzEBJwO9kwjWJs+6zfDATk2quEFhltbrg7pugF2BOZlcq+Ryf1b
5XvX53KwrXgZOXRIzPqSEKHb9z4w+VdAmAo3x/46O/67q/Q/k8iq2gP9HkFv7njkF2sZlGoi7n9N
kn0VLwQQCY7LwYOEITl+dniMIYI41/ESr06U/3d7whKptk8jOnri0KcHL6XGRPI++ghicXy6pxTj
8cmDxD+8IhJxPG79S4RFu/8w9KWOG47jeaZFXIs9LIOfhIlNc5nC5P5Fv2J5Vb7eE/dx4UphRevI
G18fvfj/3bD5jqziwLvawEjRaKvUX+Ir1DyXJxNXLBng4ljqw/KyZVnS0HGpd+DDGSiG8UY9WxR0
kQFqEXrqxVyxdCuppgQ0N7lfjlofGWTQhI3NdmVqR+PpDtNurgl8xKPJxyC/G/g4fjdIuQEo6Dz8
T3cGx0V1q0MAkgAXB47NuS4jIMvLX/S3Tp5XNTbT9LcDcJVi3TedjWMosEBLJDl54FJrGNz80mmF
IWzHEZOXCLWGlg4jPoP4vLdzfPScO6aoS5p7vAz9MMeEltQAwAViXDmVDClyPDLoDogBdFjcfhuw
nLcaoajxDvP9oituRyAM4yROpVF+SiXg6g0Uj6kODz9SIadD9gr5F1gJu/JBM03sWZvR8l6DraQU
328wmnoZC0J2zrv4dLjfRGEoMY8bXhXEsjjFEqlFlpUSMSMBoS6oh1ZKZ1dKtklrTLVlm0epXdWj
CV38WgdvRV/nDxs5uJcgef8YdNhZpMO+aW592bI+RJo3FRR/2glSbxZE6p36hqd+kAkBfbEiiAbB
cWJwmK6GtErtM4Z7HD/RwMqQZ8yHoZdH6p8MNZtz/7057LD5nsxi8wLoBce3NYcaY01I1qtJkZYy
Qbc/hvLl5mU5vt7JjeRCKZxRakZ0s3NgKR8ptQUj8BATBpK2j/o3l8e9S0JG4A2KoqO7YTJIT0N7
jhz5Y4kzml5OPtjxD4W8hqs9XjGg76p9JxIZbV003rpHkjsXU5891MHKtTgLpszNKpXpLrD5+6yC
oIYWdD1LWESoyuNpo3dVuZ4fctSDIi4/6wvCyMbw76w1MoStIpPchxDVZh5LdEddpKb+CZES6owy
2yxCKr+sjpfFqMfX6sDXALKLZ2uxkIL72rLdfumBCoFdtT34P2u+qXeBZjtOqBkl5zZ+eHh4RMMX
J0v9kNhnALOvtCXxDy+Xn42ffd/BbJhOBihm9hv0KeuUMtzqWATgyKjRQHqbOz88zEhVmJqK+b3P
6mx5N609bL4qLcNtCqzcsNJArFqvp5PH1YCH1qTKxdG6d0fJoY6XfdkDeHkoDrn6MhFY8LULeOVj
N5qXHHDGwvhuq22AEBg76A+w1jLE7RHhctOSZs410rAWi9uOaT9RwMOyTF0rKtw/nT99FfkR2slN
Rgn4JrR+qLq3cuMdNus9HTxTKxqbcR1D/l03mJabTMVUxETBr3rQ06IOzWE8emyIwPMmPZjIFGUO
5ylC8dtzdcVhw9Wbbffahl94oKv+n1kZ6AzugbjD1SC1eo/AvPtqP4ij0asN1u7C5UsCLueuD+AO
7rJtXFLM/CoVgOGz4eDFDqGZxf4/sgmktcS9Xbo+CjWsHXXqw7J4JH/b/w2ExDklTdxHPp8XjV9T
OPz+RMhRwGFAo/ya9gYKoPHx+BRrPEQCzrfu9xWUXIaLw+aEV+yvSQ9I3UNTtiB8necpuhFnyS7J
bohX1/pGkg0uJOkq/Y6beY2E4EG3kLtql4wfHn1tp0aV5g11R4/MAv6SDsW1GV23Ti4pvDUyGokx
5L0vWPvLh1g0zXAVKNsHV0Chlo8+5JyBcUjVbA1fgf3mAUL+xa5qrzfnwQ9uwHGxq3KrEA+jF2DV
+HYMa25K9hB2eEiLhtOqYA0cd1af6ANONDmh7aDIwCDn2r+usvaQJ8NJi+Aj8f3KJ6UiaBPTy/5s
qcdG76p0RCvvPNUnASdBWyjPfyW/UWeWidC0CHKIZ2zF4A4RXQX9tZFOfmzUaZwZs2CbjDdZUN35
Eif4AbxMl+qoaXkAUvN6tX0OhBwWIFx0uYU4OUx/xnc4mj57X1hsbk+nVps72iXMc6hCx5Ve7zZ+
X6ygz7wh5bvBHdZc66UEcmff35T9/SyyR7W6TZjOR8yGvlk/jAYNLCAnWiOaRWrGDDFy+qn75VPg
7QSEZ1bxRSslr3Su7IZmys6aK0C6WVYSjKnB9x12PLeGT7/c41gS+C4UY2I3txwuoU1rKlHLT4Yy
`protect end_protected
