// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:53 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bu/FPGI1kZBoyPpTOZ+zjh/sZc3iwpWTBeZ7qJKesIbBI+2ReAn5ezfAMBccANGN
rO8KnCyegHAaenlrUASBfZlbxLiral/pYpwmTC+Jl+3aKF/lJQPORInAnpWG6U5C
kdeEqRwaQw+XpqS8AiW2h+KFGEUspP5Fah7xiUz8bZE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
hXQjTlxKDcNi1rQR1UstNmaQP7U7WsbbKlM4AR5vFE2iv+OUj0mZ+7XprwwPQhVM
8q3ywtHdmaNPAeR/hdq8JVYwDLkB+5wz7wpLh8gWCMgII9VcuyP62oOpyj3hQMoL
1zxJwfnUj2mj+7s6U/DziiJcQcZPAe/1iyGFJrYwhUUBcHGwK/OZLGYTMcoDMP4h
ax1pYs8sthw1k6T3ioD3sUkADNzu7L0f5h6NihAavs1v0Xs+QpWpxDsgieUjjThK
Mshxc65K8AnvMf520JraILMnhbEKhAX4XyHqWrXyiNZd4pKSCYFjn5miD0Rb+kYj
lvuW+BYluXRJMAiAJZLXZQWxtWr3byMQDDyBh1eVmg6S6J3dnKG05oLmncTNOqeX
nSIioT2oojXHimRzpZQr1yE60uab75PTCkt42bh043ozHkp/NNO5EUOgan0haWJX
cMDN94EAefOoJvBc51ItX/kiRv5+JrAWuZgLwO/wkErDCAyxVV8H36Ht2nq3N3T7
lgtP2CXe7/Btj5l1GJFXtWXgDrHlYQNSZ2UsnNmH8impZYUSJWj5lfF1/49s3Hs2
6j2MwZjZIEGEjD4vPv8xAHuj3imCi01v2eR7c206AHhzRtvSIVoJv2DZwg23B1qg
EJfTxjBOUcpWwpCoBbweZlMzdeX5Ddkuhd7zI4/Ufcmg5WCXA3WiOPuArxZKLMm6
+Cg/ciC4rsggJ+6ADNJPm4SNbrR8yHYp2g5X1f5qjUWwbWOWTNXCNxJA1cq6PL1p
wOWEspuiyJAR3c8Z9Vk2vKWQRxxYld/Ae8iZORQkjVVaR5awE25SnX0j6eAsd51S
I1sngWr604dK9KtvvsjoZSvw7kZbS4pncr2ImUPJo+NCFISFkBlUAtDyE35iBBfl
KyIPR0blmaUqNGZc83RphDCWspPcV9tuWk9WbKh/ostC3NAZ3xXVrrD2baqjR4hU
tm63NI2MFcVGU0hiGyfHGk4QjUFkfv/cns2rPeNBhOUA1a/42N/cYvNBx98bU5AY
ox95yOuRWh4DcC2p0SS1t4JDWnd7zY7iq9fBwJho504Y07odeIcd14xBURH7HW13
jM3OuyPwqz0EpZl0A7YoO++Nv9hF8StZdydM6w2BVuubofFvPl7bURzznATFm0Av
7bBGIFjDheOWgEvxhDmcdyKS13DenZKK3+gP8riZ5vSi/Q+yUpjn0gwPLXYiozYv
ZvvHIVj7q6OGzkQhRpH+TJr7LLy97ac+IsDrqrn5cikXOwdzmJQGUYJZBpLEJrM6
IMKKVrskNbOpy5ypAP9Heb519GwByUhwHUbZptfZHT0H4n7QCWzSrYOy9g9qu+Lr
f1SFv8zTpD+wscXAraYvDCakYUdnOXgEELxVtAep/tu8svxXlm3Ld2a3Dw2Gnc8j
4Gi4K6nqRP3wChwVLtZWfYIKIUx5/7Kh/NuPBlUqehnP6pUujvP5Yx99M77JVbkU
zWqMHYC78+IrXv37F/sGqSZMqLPqWin9GwSTsAHb9eLDAgJe4nDclmEdcekwqlfX
Npz/9zmopsRzOkFFP3ZWz2EwYqIDCH6BK5tjjeNZ3U67DuH0uIou36g6VNo1cUXK
NbFiuBOvH8Ov6LOc0bW4FJUZAClQeyCR5A8GP65mt1cnnxeIKA2rFzMJr0Bs9k5b
mmqzy8Jh2xWuZMX/FkwD3cWfd59uv18d9CB0jmDKH99nIshCgOj4DImnR6kEYxwZ
vYznVGdv+bRGYGuRqftjU08BvW9XMjUNbzKTqIJeGkAgBXDrhyRRSFVGQ4KSy4I+
XcQ+1PreQvOiRmP582ELe0zY6rHus0OJ3su1ffhp1NAtQQm6tTCjVbHQq7sYbr62
XpjVEnMQzihmn+5vRGtguqhyAfjjGBTf0wbCF9QJ/9Zq8DUT1hkM1vZubw4+OrW6
nXz+GQCcXG1AOpUv55qNVir/PHnQtRprID+80SPfRNruHA6saUuRdG/dFWbqp98D
nP48zJZUa3eIvo1wQ46cTEEnqxyoMgj0PJoCXSIWQPILS7SkA9C0uPjvUe3ucU61
5Ok9WmmDcfvEmKiy8pf+1Grb4Wo7P1Uw09VUSrEFdFU0+jeRnHmCkmQUyGLrR38G
2e8H5EILSFx6oIHH5uEK2dlhIk2YnBbRn6DVwuKzcWjhpMxLml8S3gOOXAlP+CXQ
iJSh/1Hqgqfu9BGwnnKS5qIygc5eGx6i+mQ2/yM0I6+TqoEXYvuojo+8H4Rt46JI
7NnFFYoyap1W2Z3ogMalFmqbOhFDvoRC8DRUXkmFy0k7YOp53NejiMlzQoRT1uhp
DPp3mS9oVUoBkFHgqP5sBYWz5ZpRoBwHxkYgB8mYI8GvDh2kmcqG1JElX+TCse4y
3ame2XBmaYSscMDFf0WX8/sByiHI6+EHJ13BCznFsZ9L/wW+uUh6QTQvrAiJ0L6X
ZT67ewPfmQEe2bDuaVcHeWIOpMlKaSt4Ki35DhnBUw2Gyf5IQxFpdeyFjbagNnck
CC7V6wd3zzbmdHawITy++KNgpZ7k2m3B3l678zpf3nt/cj4ZqasJPUpqTVqMSzLw
8caMo5ZbSUTx/fH5Uk5FgIMbMY2kZKCui4fP9b3YEqsYiBD+7FQj16zCQZZRh+YI
QD5W2r435SukCzCJ+Zlm4A23dV4D/9QxjdFIHQRQHzVSsh2E8ia/XDivO/QbQ5S6
PBADKr+O3JYEyND2fkfpic9uV96K9tT9qfoOa2XKrpCg+AT/iX9wHPkCltmyWz6H
wWVnEE2LvWQLEZiJPURrokz5btugUQqxu2HS/kznXDBXGK5VhuuVMjxcQXz794yt
5FL0/TZZasHnBcJBDcVBScxJxhYPZMGF4ONmXXczPLwnpqwpZiP3j7ag7fsqRkUu
cw+YghrGf/awjPFAmcHdnmYDJsjTmiLD6bM3cJ+ry9AZr7YhDzc/0TIxyRMTJarq
o9Kp32dFH2r9VprJzB4Hr1ztfPA+Z7KK7uCtOnywioprCq4eVLtOZi/mREsVS3lh
48NnaLi/t/CdAs/Vo5gguggpcm5EXoEWJ2orPbblqg/KuchTJgPWpAklL2bI/nUM
NpmmuoJi5s/4+Rb3+fluHxJRGMRlLzg24VK+fnb4NXyWdHjm8hzPEG+LJ2fFx4DB
v6mq+9qtUm4pzj7LQkkhs/JG48rW0OY+LbP0vooXovoxcTa9TT97dUtbY0lPdWyk
eGkax6HjfeGXbeSBera0kMlhrqBw7FEgH2sC2CBUc98Wdd0hUw4tlFb376eeSFhf
egwfh1ZzUjaQcMs+3yJ86MyGAhl8nsz/LovirjlpwML/H0TKFuDewniPYfqTwUqJ
8OR55JNAWY/7RTo9mKqx7Z8gL46tJzZH2MQ1JMETC1IN+25rIHAj2/4jtyyKdQAt
GiEj3jK5n+PZIQ6jNg8mKdRIJ9Ttil3whrcVQjlpZnEvuJw3xkxe1AigSysSXRg+
0ds5ZbR6sRD8p1d4cooDTWB5mbAkF6FfezBGnPbtopengn/zD2jdMXQZgMUkKH9d
vXrOuDbIZ2PK5I60dTRGY2zKvPWNjFaBkr/LaWyiwZr1/kkXAy2yJzfnGmpZRuBD
UyOmNjyKQOYaIdvyCxUt37eZi8BinaTYj38j9xL1oUnl/xxjRMPtH0KTo6t2zEcp
i7X4t1m2dx42F4EeHHlNgjk/Jhe0gNtzBbT943LN5wzr/dJPUwoFLp3VVuvDIlM8
pXTYdQgSrho5PwsY+mQKhHCtXzgg825KrjAWD2+M6fj+au/zGaQBJosdGCeQa5Fy
X5On6XH5AHRfGBTrBidWEQNY9lgf/k4iJXbYWXUdTO4WqgPLYdQnWBF0SmGaEfxk
vBc3gIC2anhLzU7GIdxIx2e4myyBt2BFPLaOT7V3mQue8DyT4amC9q6SXupjHiFQ
PRvBqoGgtwESact4Hx32ucFVwrAZgrepw3pwRR3Grk6K2CNR8Qc9IsqD3WPZQM7X
zUGVHemxOwE2UyvYcPm2xIKnh0bWiDMbPUQhxXRUBhNt41UxuP1E3kipdYo/rmPY
WLyv8ikVkSbzHiNv27Wuvc1JvpBF0PedBYZ9pZIpIf4Q9xrUw7/BnH6+xd20wrgB
hIKrfkwP5AqXU9Xb0OU0ku78bFAEmaJ/Z2rWe4U0tFW3BcsY4lUtaLyWlNptfSbK
DP+RdUkp3TpYZ6X+/fkTvf8yY95EK3SJS29uDp2lABlMeD/Kb1zeo10AZbQRl4s4
7jTfp8ed6/6whHMgIRXaShP8YX/fPXbuVkRiHoADJAlr3/08rvfnQgly0fIH3SVS
O/3DTmXuUJbfqpPtLnjNKWZJiH3g/2K3kpDG6XPlBGbaAteEr8vqk8r1d+k6H4oc
t8LdBIBFAhuAshIFAN6rmRkAtp1YctMBwtA0omneJJlopo31W9zOhLKWd9iQGBYF
qKJWg74eYA9mYkpyQK71YuKD1/7lGSTFp2wziPtTlqwZNIRTR5+kaJMa0FgpATmT
jJb9KfIkWK7qiNZwqUjjZy8lqKKYFIwtmhwGPu+qRxgMOTmLrELGLOMd3UoYS8Zs
3RyyvFxjUdPEQmGwQi6uFaaN4OQ4ww509i0eSQoVPA8fCQim/yQKqKnqboyWrosg
pQODOwKR1oAJihUxbW9NDmaejskis5+zmoSce66BlevvWEAOgJSFxEGLxQyhRQ1n
oR3IwvvNqBhvNPt5mxc0Izw+ZwpXjRSx4ezXu0udtsOnmmrE/L7+19eypo/S9kIg
JVRHftg+tf/rJfBqXOr0glINVC8UURCwP/wArnMFKT0vAgzTDMdylgbewuV7vHYY
jhyyubqZImxAhycjXshPLn/8lVDxFHS/8qDVEnqglkIgc+yQW99b6Um6d+dD1EoP
dqxsPxUu+zzSVTpI1bavxMkytBaqgRQcTrClsBcO2LI1NzfD4rDkTwMy1rt2551W
9FRmT756cjPViflyCyZAv2tEBVz7Xxcglv/h2g8AlP9IShrbimKkiphS46xwIRrr
CDuqn8PBhA/NjGkO+6/+NVswfBrnz0nijxWlJFxGgmi4ohI5Ug4EnmyNL52GvNdC
MF5AtI5T/rAhv1wYaDxK7Veglulru0Y3X96bUZ5LO8vcQPc2c/hs7HFUspEa7YD/
DriNsLr4IbhOO9DkWewdfa/zHb2neqtEzGasK6Mrrxu3DBClVNZXKZrR9zdWH+qY
AWtz6hU7OZvjcpk/mT5fGhzK3nA7D+9IXh39TInSepmCpy0srCPPDTEBcmvQ9cqN
VNua/f73dlIRvsrMMZSwXebYRdK1/81iFSmxHVaRLQp6HmecgiXx5cl0UoY4jWet
uXR9UtumtX2bUrcySv9pylYkXgSeyJU2ALCJsmHWDo+rBRzxZTapw+EpdsWousaM
ZIj0EETWcPsAQ6Ub9syyoLosXXtBZkJcA0QfUUaOP920XKY8QlsBESU08lkB5+hH
Ox2Fjne88FnpJ1iyHJ8ZfW804TUclqSWDbWqCXdwEsYknlgMBNPHV+ssctem+Bkl
OSyiU/HoTzHoihsSB0UP2Dh4Kv857q+tsY1cxJ0/NcG1Pr1Jc+vCzJQhUG1HMVVe
i5niRQyMb+aPv6l3vkFvKhbMZwk6WXtStLDbRNi7bWLDw4fo7nBjAnKJIeYpc1Pm
TU1xx0roohWWigViczLxj0PDetWedgUvhW4SEWghHZ/FVvdZZwwgWVDwBwXwZZMl
zzROV5NGnO7mCbAzq3k2B6qVQVCBHZwvr2od4FMA8egE1Gxq1TTSEz5OBp2wFvur
l0aWhv/mdUx8r55xOEyOrGqt67VMpupL0Uo/oihJEi22lymK1UeLFk1SccybNj5E
EyiG62x8CwVI2d8opOk1iUAQra4cWNl40qZVg5KS3aBuBYK7nWU/wZ+O+QBzCIxe
+DRkB7OA2p3Bhl8ArAFHSy5iwu36eOy06F+6joP8i0Kp02xkVnmSzPs0z1ARh6lT
2ii9axn+/GjckRnFvVJLhu9jcWn199c74PejwF/ugbQqDyAsP6uPapwGLL4GvZ54
YTQ4td4jb0xWkSZg+MXQgfYFlymQqiuH09Jdc71/I4aDQe2uF9DcXHQkqpMBoEB9
0irm3CcuRaZ39F8ThZjE6ieO9fNtjGzYOoJQGeNyxHpNz0qYg+L67ObPA6qBXuxq
Z2lyV+xBykfvlIW8N28ps2r3ulv07/PXEi50LEujCHXvGDen+olhDlMcF8iOTMOg
YxeASWFfDyKRGdSdKr9trTFVoi9vC9+o0e19086TkUP/+yD32K6ZX5aFh1N+bL88
GHnwxA5AOvs6I8LG6qg7j8SFdx0SlKbZrq4KM5UNRTqh4nF7Y1Uo6bZJyVaFyyks
3cYNZx7UQXPdaXs71KAx3maStjKKdhfMnttvr+tE5agFQb377WfjzbtgTzeMEklC
Kmta8nI+VBrJyR33k18UL3jYecaEQ3YAKIz0kJtU9FGuvEwBam0F2P8AQDqcMnd1
Pzc2pWCabx+UU8MKHJawx5sofWyO7uRbeBkVdYyoDuISQ/ZPLrLptf6ekG8XCWF/
yAzQPE4DZBAoPi4Et2CHgHeUsLURH0SsTc1CQPg5GU6ibJ7qqPZZwRsC1Icwfsmp
X9TnEJDrsWTLl33oZKOq8893Dyvdf1v8QrvGqyLKgQlL5wTjVyK6Vn+U+wq5lBVw
Qh/Oxzh9eMvwysMFoC+5LrqPLSHOfzEDEIN6Jij5Cd6qQumEmy4n7F2acVVW0QX6
mxjSeM254Iy0vZ4M2vDxIVLKcf0uwhRskH+aGjIR7TELSE8GLz5a/NtKdsCol1+4
KMSed1icafUReROPL8dzEhd+fJu8ydAtxKVXk787Cqp3PhYiIU8UhYWkmYIcIEXE
EfXVQseWgp2YxfoANMPmeXS9zYF07C20paA20Kcl9yq0R++weBW7RuvQCJxd7R1u
858ksDh7Rjy5G4ffQ5AzoPgPA/pVuhasX0e5LN7zIuUBU4cm7U3OVMWjzxcElg9H
sfKyrTAGvJkLppdsWg+WPuHJ1svswzhu7xrOAKup3JH/PjwDrzyxwNlI9VJu56Qn
ECiKnToAKZwi2zKv2pcvhAxXc0qlZ7ZMHOiqFTeDqfOyKj5xM8I869Xp1erINNsq
7bHJ58+lm95xlCNona6RSueJowP063dL7uxUpXtQ6W/yaGJyvJHi+Lj4OaM3XRUt
y0SlAml6l1NsdJ0fQDUZljT0fYyS1YGyLlW71yNI68z4gz8m41QI9jkcgI9KQseV
85l5GSlUsNfIVpC8S1hCDAfECuikhoXF8R2F2OeoFHBjaSv7GrbRFh4VYDg7J5Se
7oTfV5e0SAXYalLQ2gkM7pubJRBJ+0/cSy1+n6kry9YQNbtdX8t4XVqFxOrvzwpZ
0q4+DC5BkbuOgK9Ac/Tr7wB0o7G8e6tOREIlIln0l/oIko/ZMfcWd7i5aDlVBwU5
WqH4yojc0CQt287ZTqjzfZM953JvWJbuNXyrgGk7aiiqzZ89rkGPXpSfn+yH5hTS
WDUYc4cRWO2sYzkENvsr0RuJMmhC/pUKkVqT72A5WbwdHaJVVmm26RBog7uiq+8/
EA0PAAw7i4ocJUBWVtqY/YclfHFQXdhe+k9O5M0zGwkPYsBispaNzbVcVxWbkukK
nusoaZ3JrXCI3g10eTp0LVtR6nhb6Aa7sqfjqPhyyxK6/geLQMq0I59y6mSY4j+B
n9ZazYmUgnTsK0fqsM5yrDyfgXqr/U3VOAb2AtDFIt2yhb8MuFZC0t+BliSZEyFm
h2Kvi4MvMeyDjO7Ug+thaChLf8dVYkTrembSjMF4wyg3qhHsNY4w0sf07pVJ0l/u
R/26PfqebXYIx/5uWdjn5JSXWDomwvfS1eXgZ3hnJlkmavCRuRiPFqHn/16oRG46
7F7vTb6sQkxBr1MPT5EzKOYptN9lsSk6AKlC9gRbjqkN0pd7ySCTXDSsGjL1SrnL
VE9A17XBPVNjp7UvszrDCxHNROWYg2i/wspu2yDZxvZkwSVspGHXaMsrp0hKvNfU
OBetz4Sac+KkKvQIvGOaIvvroegKDYxWprYiCcG7XwyO/RF1UOlKgYxAbWXV63QM
IaJr0jdt+FrrwbHi8w5GvPMAqrme8ouVkH7vdoJxp/qOyPi9wBwAR9+xGB6PaX4L
uhkQMQePS1lAjmeAIluYRuJ/qZbrupjjBPd6jpLSy7y3Sq9nD06xOzyDANyXvZYK
/ck1B/l0ujgwiCN4UP3PeWdearRX+HeZ3/kfEc/kkdJ3tE/M1R40wxvF6e/WpgGd
6zDtjKFlI4FofrCpGKnGS/GxjXEJpzylXnZsdEhkyx2fXqJXYavyT9a+0KprsAVE
VRo+npbIRZzaAyl901WrCmkr3YynWLJIGtpmJGI9uNyU1BHNqUUugqWX2ZxaYlrO
bhaGAbCeQeusPTw9+oZMXxJxiljt5mDPdTcLP+zZxc2wtHfSq8yPSdUFUey6PTSp
EUX7TnXL1TBjwYvyV+5IIMLuWVrfoDbMIjWYFmAE1ZXD3D31NHbqiULdW+zNI9Fg
ob3B2W1E7O9kvTKMTld4kPN5csQZzwc7ygczcEUw4WMoDj+UFqRlIUZvQCZPtMOw
Tnkuft2KsR0qLKiz5lBG3ioFxnfr9DOjm481AbdB2vUrA0iVXN/GXbldA2fzXiHz
kEf6Kagpfp6LiR3a1YelzHCP2CbfcmCK+oJrfx1jS71VHZjgs7WSzDvs/FvN3RJX
EM6Xlqa3VNF7sZkGhq1kW05BKjkWcplnx1re5g4PtdRpXHJaWNPNd/TuvxdMEUri
C+QgZ7+xJsGTjebmoa2NXgX2PMLhyM2IxR/H3uVInXivIHtD4STYVG8rVmIbekkD
Ycfw9vWae9gkEwrcKOUnL5pend4t/mwaREy93oLvcvtuZIDUt6TkIrdhNsmiQabE
sgaLJz9K233Bs9WlRcvPhPWz1yYjYm3OWKmp9V0xxuA7uvztLtp85RvjrpqdNC78
WNQvLVSLrpsLD/S+8SMqmWEy+6wY3Kq2qL7CvXak9CLF+CdHGih08LN3YDmB+XYf
DscBoTQO9057+0rn/lwoCfT+vWqL+w5He+w5ixlfYZBNIRvOPkAt1FwewPZIEbMe
2xwVHCkU+PrHT9amGN5JrxwWfZAyHFII1Rqa/px335L4hf97KFCvqtFPr5iP348f
j8K2oaihdUrlwj1afTYUVtJxGKWPutjdoW+7W6Hi0DmQAfS4uX6yhkmMd16WGewr
nP5By2TLMB9bL0o3Cx90IdPoJ6W2CO48EOdn+pJ8OKZXHQCzEVHTwTo8jV9NCe25
TyZv7lT1C9KQz3iGoClq5xo0wIv3CVZiohd1v3JoSiB+/1d/0rfsEHR428b5fdP+
NgzfYhCul6cHZvpmK2u8H0pj3Mdo7Kn1huXZ5cPA3P4wdoWCtUIipZLaf1uJOe8c
V0G9YIus4Z5LCvEnnA7I+NW3WPqtRjK298vIiKK/m0BP0WNJV8+xpV1jQwgbV+kK
hLNIbqdsjmQlgNCscGKUGcB7LiY+8Ur83d4vE+V8r8kRF1Fd8FLplwdt/XzwKg+0
w3XM9hYurHL9Uaj1uoPxBGpJdWMGSYCJFhPhLr6b9fSsRirczPSrMB9lETtnCXwY
tM4kwDdkaRSyAHuMXg/QcF6NURxh9S71ydgNlGOXXLIj8bhuchB3ZZ5eTAAFUjNe
3GfIT3vxPrDb/DGbz7hC5SHegxJrGHOl/D0+/AVXN8HblSdpNCbZU9yWWiKojyZ5
Ckm5lx6eskjYAq+u7t3lMw3vvU1Ih9oPMru84TXqy/Oo9GWD0Buen8QY5OxOgjjf
N7eslySqrhb1tmQulnJ59O+ZTRrueyVREnlanty6opEvjpuTnRDiAERhSYDrbljN
5zMhhrv3YXUTc3ArnUbs0n9B+331ndG5xBynQFI1lwDFQeePJmY1QFSt3JpiMWGY
IpNjFWAurqoqbeQacmGqvF/HxKS68ehWtHkD+Ilx7NzEorbCgYNdE+UDWRZ33BaN
B/M3fdyeYoHaLROkb84Z2/H7942wozisUSYBXRzpYHJvabGy0EY0eI82RSnALV9y
pqaQ0fJ11tQJRnNU4oNVZ52mpCYBN5j4gWrJb02hWwQJqsYnRhMpsP9uXtl7Ntpd
dBu/6ik0Iskw3dxBO+vWsuPzVJ2Usf9d+/Tmolv9yX1kFiugsTKeQbNDBR6prZ3q
PuGVMn9MrjejayQ4OdXfWTv+4CFjSqIsYFKn4XG7L1V8UzzpEfbL3CTpA9c8VttX
PoajCwQnkitNesVTAhV18ECLXM1VpBPJ+VdmBNUzROOvXHOnOMkq9p3BJ2YiGB9m
f76xmcj5Ew6Uk+j3vI4yZ4h/z3qpaclEgg+B8/GwZmvWKv158XA0rnS6M3ppPKTv
+KMNT4CGQhimZmDYLOisT3N5jX8Wgq4eMCyLRhUwQVZRNrtRS81l+MvL9noVVNqN
ggA+cxxYEe/3ITjt2ROidCOV5PibHdvaWWM/qjDWRRQOdqrbHRJ5y/XcHaQse1MD
uEoQzY2+5mHwRXg6E5wOOKjmomoZQsJRJ1wGkrKX9wMx4qjOcHAK31OQ5sKZBF1c
LlxC1UCo6GavRfeDhzglQAjxX4HRdNjGVxfFVxGkBbkbdw6JSoroiaNlREIGXsJd
Cg5RuOsuVPpdUTWK5PN7wxkmDdXZdlH4h/uVrjM0vrD9dK2X8thi7mwgKEMa/SAb
GcjBvJtCae9QZ04bG28iEM2BCuVPk8lkvPsRrMIYAUQzxoBitEu0BR2BDLUSsv9C
RX83g0X0/rfneohxC5LZym5GCWMGwXiYsnrbOPQIUQdiVBRTXU9mT6/oKjEMzLSF
5QX0UpaOhailS7+EJspo65g24+iNmrhFJtV3XMalsVUXMmKCV05im4p41RTuI6rM
5E7oXpvKITky1/TXTYlotZXz2HttnuEhHueDEj2JpQmjnTbesCYDmUT8ogj1vdbZ
JWFAfxdxuISoS523UDqpXKbxhf+UOVGgj1oeYIh+b2qo+idKC3SDhMt1obkiJAEf
NqsJ0BemrgnN20CMMK8bvK5EqvBDFcvh3JHlMkBNEeA+mFQRnGRFwg5KOdQgWtLD
QyzIoH2rbjeH8SDt/MReJIeO0msdmhPFn2dD4AHQ6ZqOLa1JN7MN5zwvtluaDBZV
sNtXaORXGAbEvQOiphl40gfnhj0C+3ztqd7GNDTce4p2IqcKcPcSddAnBzZnFRz7
u180BCh/SkSdhY0HWUbEXxoerbycPZI+jWbvb2ZluWN8ru7YehfWOxfBT+EEszOt
RjODVIsQYtNFmgttOIws1VMAECjXBXDLdmiCq7iQ5L1tmEWlM8F8DkbjME3v0HXc
jFnlRn2c8tZ3ba8jnGNoV3RAQHzJosBG5HvIUvDoxbn3tt0b63knMt+Tk0bh69NR
hb3oJjlnGBOgqTR2HWAz3FHRmCFwOBcFISgy45gp4Wivcz5smrj4GJP+DpQNrRy1
SZvpjGdzLZczxAYmPv0hKJRoW31+TGWgcbA/MZhLAW6gCgubzZ8gDvXUFlERlkma
c0cTjv4fjuV4GW9DJbflbat4w8DEkKaqSDpeR6eauyuZrHQFBVjDbJTfiIYGK4Vg
yGHYmtkIekdpvwZrruXVgrUKopny2NfPoY95sXohs+zSYB4OrmZFOjmMoPIO2WBh
pD+zvBk8uYXHozL0dmKeiMpNHglzWVE0h23DcaZmPOTddDd6WLpNmCzD0e+INuDY
5gQDn+kqoun/vj69PJOyE3BzAt52gNTizAv1TFrQgYN5Ulfp3eG1JOuIn4Ez5f6u
9CvSEnw1s69Beldt+7ZRtx9pKo7IlAJN8727pP9+tmZj+hJ0urRsZPs4KBYd9iQ+
Z8HR2G2TslKuGZB1lveK85clvUUS0xvTNApLXktA4fcCvYOlAOrj1RYPiPiglAQ3
OSw86Tc+VR8vf8escEu+fUCK1Jyrpa/QU/zcq1rjZtFHI+re5wgBhZoRXl9yKv6O
0rU9uCfXvkU91LZchIEeEh3pHIK7N05T1AVyNHGRiMM3LCZufNtYvgu90837mjkg
M/4Ezir/4HOyVlqDozyrz45Cvg5vrF7vQb8QVnliicAyIHKroHMVmwvRfS7D3a/y
XpUCWNlUTnPN4zwJVh+8vg==
`pragma protect end_protected
