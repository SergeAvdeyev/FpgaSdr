// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
OrMHYiFRKQH+T+qUKvEttaGpKj8cTWScC4VEGRgd2UVB9ihJjzAkXBcMqV/ZukhPuSOP9L8gxJtU
fp1FTRhd+FuZURcAPicPnJCtzLAARSH2JNOAUzledB+J1NCd++7Tx+gknwi9bC4DaUaAdOadH+Fy
Vsi72HmgwZh0Iz9/HlkzLaQNTdeR87L8cdgqfD8svZ5+EHB+IAj0yxliSv4REl9Y8mJnWKNQGYqe
ZBzoY9Nrgr7Hlom/vrvdG/Vx9K2W3NxjTeWYT3EptQBkO2tpxqH0uVKt+sOAY3FxAz80OyyPiIm7
Rw9qPgWd0xLvOv6t6tNX2+xm1T+SEGNrAnx7UQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2960)
cXYFyR//OfSXV8Nzdq+to3tLJZxt18NCbdfN2CTobBigS41SPrHfzviGsMjfNWwBBN+8FgWmpSjd
MFQ5n4lzbRpJMGx6Khtpn4LKFNn4tMPUAZc8d4NuLsJUDWwWJUb9rTBBH7cdiMdh6t6qedZztyi3
Zl3z5HqRHgwEP0QJlHBP9UQ2oqO5Ouz2BjU8ZufCiiUhfRE+PSwNXaeP1g2aLH30pqVwz0HunkER
8RB3XPNV1oeNzMis6WJ1TfhKv8gN3O+UNA3gon70hzfxs/kJBvsRvxChC0zjlL0Iid8/2kd2do0v
i7oclfmzJvUVCfBdXo7iSOC1+Vrl05N3CG+f99iDJKgNCQEpPUQW02qUfP06pvHgYB9vSMoOEeEV
yVUMxCCobAUtR/1xsPK+1DkvvN3lyOFBqdCR+TNWxBH5L2UUWNpRvhxKCWQXVUDKJRyPhidy120a
U3tysOUJIBpxynjwlP+zRJG4MbrloQ3e08A/ly4quYiMUPGU0ifdn+Ol8ec26oJB+4VoE25pBhSP
0oCHYX4FTZQuZxiojhQdmuPECOE+lmiLnGNmEhjPOYIWvA93DLNo3ljw0PT+XY8O2Sbik77Uv71f
o0ZFnFSdqo01JLXcLaWGhKXRRDoSFnGDW8H7Oj78noOa0s9pRDDBjXp/MAQDmkzxeDNWeIjtwqxs
uz76l46c+Eqc/82fOteszMvX8pydoWGnaYsrajZRl+9CpePfW8wuEe7DIE4mjz+V4Basd49W1R4D
OHawXe4OiskudznDgumx5zXFVYSVu4oSPJzhD7WRYiA+AhPtQeq2FqGyZAwROLBxJu5avF/vHvfC
0L8pxpOG98B/xfPKTpjxptAAC8J0vgk8CarJIqt+5cYFnvGznOLFKW/tq78j1w8Aygq6vcfdWmlw
frEbGcr/wqc/PThqZdGXph+sxcjcUnrL6INvFKZRv+9KLXUXDhSBATkLwNQ3uRe4pqpha3T0FY/W
7143MguJQeeDhBuYgeViCP1ZToDC75U65IGq4QoxgZNah96kWmkRk+IJBJSMonMe/gohN88dKRb1
l3RZUshpod3fDXiSMcQW/GzQk7PmEPisnY4pZIsXy7UCleZcb5MVAb9DB2dCca7Buj81Gsa+UNoz
hdDgLxXQLvvPUjDj6WLE3S31H3GOp5O35bMtnzsNF69NvM2g2jGvmO11DfNKSchb2gBvWLg1DCUW
R3/rk5XNjdD0a/mWlo0dJH8I744uKId5cjqOn2X/opK7Fg/9cgyE9bxe+uG3U15gzMmvcbQE3Jil
CrLe+MI5M3ctU6ehEsBak42mqF/NdjmxXIxfG48y7WiRteIG5gR2rh0/BRWM1eV0eUNEOQxoy9d8
PEcSdNfvcNVffjLDpLGlhtKiA2yYsMhFhMo6luyVEvxpETEwLWgp8vY36KI8S6m3Pm4B1H1/6d7/
wRyx4wXWtC95uWclkc7zJIydqylL2vvOP4jTuS5BrIYHJfSJ0cUnauAIzX4LiI6nuzrF1pNj6pFz
ZZmrQaHRwZDfHOSsDcLneCMdzygLXGbMKMG6k7a3zbFk4KO3miqwWnt5jhX9zQ53v0Xd8Qx5/2yf
ZHPbUjrzTILb5DV6Z/ItaTqMcE3CzcmJCmUlNV/mnzXBr//DkuTH7YCMULWTafTUF0kFNd8Cy1xF
Y3kbBC8z7vTeXmcp3+RQ46mQO5NDH3Q71fpedxAG+OzgcF012104xiLmBAQnGz3NwNBqKjqXfbt1
+TlBS8/bgTVa3ptGyz9fNXuEMzq+LJkBmPgMAeD//Uc7edmUpNcjSj378zS4SxX2HmgePaMmtLXY
SYYBPKnykq2q9uNCQIm+313/4vPqU/9kosvA3MA0eYonhqd6DHBOSd8lQAENZ93S2HcA39BqcR9E
4vTfXIEHMe/pt6wdoQV5nj1R3ryNQ532Eg1v6US7NHHLv0VimOUrgYa+QUqhPTawcCYtrrgvZ4Bn
KYUKAe+cjY1YRJI4IIqAvqi8PfBu+Tpw+SPCoajsi6W5QdC9EhvdOfJ3eF5w6Hs5ZlOO4HtOY2un
pKE4q3HgCb/dhI8Is+CycG9VFgqhgm2HTZk8lv4TY2hzH8iKzvpT/IploTpfUXex3vAjMH65JWuN
KyBqoZvfo956wxmf8jflWxiAI5eQm/VdZtJs8LWwZ7Pa4rD1In3UDjxqDZ8VI5TP9edy1eoqCOpq
QVKc1LeV7kwpuXWlARTplCetlBcaCvweV3ppODrIccE/PHThSMeq3Dz7Zm0d2yaKwz8KyJMQB2Im
Vv95KSX7Uw1ngdQmC2FJGNGoaLPaj6E3Nbf0zMN4CUUWTcevJUvYMwdyizpqj6jtpEwKUTHWbEYm
Y4XNMgLdo4kMkPOG+808eymBvXqmagLLITCt0/GoKlFFd790q296Vh+D1s0rM16plefjyaDJcvZt
1g8WJMRy707Rct6lHq8XcaBOVdFQAA66FzNGzC5A0iAOBUjQX5KQ6VYYxzerk+aGxYjnLTjGBFFu
hrxco+ylITBu7kGx3bTGq7Z9uKzUPkQBwkiVxkMoZvGXNyR6GWUHknDiD4GgJpGxQ1eNmrN61150
rN+V/uZjzZVWKrXlctUnQAC5Ulp5rHUFWbUTmN7A/6+y2cXKrk+Jm90GqUVjRkUUZn7/zirT6g3R
oeL3EWnZmdO0PskE5knvXtq+7MjXx9xmbr41azQaRdC6vaFUig0SN+YNYUQPmOukUQCETaA9nxaJ
TaF7+Hbb1qcYNghxT8NrqzEJw5UsRSerxONR+2Pyt5yjzMk0fviJOTQbeR9/GflZbt8ICjOM/RAn
KErdG0VQPVaJB51wwansAdrhqpB2fOXAgQ6ayDHxaSVxKNO+VbTleBK6o+1zNEaYChJZBEP3nQVp
LAqgnW5YE7ijyHWhQMZ7NQZgapLMWbkZhSO+y3VDQrtAKZs5Et3FSQd8AQUJBZiSfiNoQYPQQG/u
asHG1OBoHzxax2scsSHmwzyo0pIijdx1270GYwnx3YSlxWPTUuup3Yblv7sx3l5kgClShUBMrYwK
wyzikJbYAwzAo8+YTTlTxhfsniSrn0f5VtKPuCqoFOcYVLUMHfM78AWK6DW1GCC7c1pM7w8EV/iC
hx0DkX4J/Gn/78zwpl62CfDdXjA9r+y34a5UGfD7wLUCoIMDnTuyFUlpftJyvjJZ8O9ReDsAM8GJ
Hib6B2aaLZPNatoEdKOjoVWcSzLu0LJ+wtoSkFHCMk55PZQ6gZOGDjooPPjVrNVdrrOGt1yzn9Eb
Lz48/ZkZda3ph2Bc6xBQ0pRXJ69C1V9u1zuEPb5bEEaTBxYs7XwQ4ysuBjcMHxaNjxz+UuLjFTif
bFerFYZhW4mUM+Mq+seUecVtgI89TRPbep3jW9FDYIqQg8Ia5oylFKzW0CidgWoDcHXVoMRim/Ao
Bh4IJdZ+Iq8F/KKOY9qD3XqtT7A8z5qgeWmfarDO5b9OTRkfvhQT5YeIhEPnE0v3/62+GOES/hb8
2qu4jZWqDbIVVJtY9YjkBm4zzzU51HoEcHWlUgzVkTmXmMq8M979OArpkpEB6EKw3oxQEAiJZmmb
qIeOnw6Iw/a4lAao6wMpKvlaqC7l43MEMx+Yvg7DnYKb1vceaDAPAp6Kxa5pJReXsklWWF8dp6GE
y77Zoo6uPuw7Y7pznODPqtUHTe9svh3nLHgNj9s6OwccowDxhJHCM/x3mDhl3aAGaU0F1VexhJ40
fAbRDtt/sN1dj85/ryLfxFCf9mNVP4mcMLt0cipUEFfE/vIwri0Vj2/Vx8d3w1HMv5qAElz9ZK7+
jzV3+oOLlUQSzaSb7xk11FXk9+tAkeJi9svBhT7uW94RNviM/3zP0Oo/4FebWSVWYGOa98+1Rpa9
SnkwOPBd1wFIdeyAj7+WYY0M7Giu6qtJwi38Bob3IVXBY3oR/PTkimzBIbeebiG6KzKGw3k=
`pragma protect end_protected
