// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cF0xa6lhjwM4AfQY48WUT+yEHFnjIk2a8kYJWGPLOr+3UXqFfnIgmspX3G/K+eQS
VDkjCUMawWGnXMIwKBorL2Jto67cClwyr9OxjvJt9MPRO+1MObyKoSx9OjnPFWwy
bM/pQh53YOtPAXfQbKkJ728GicIJ5ruqLZvE7P4hkLA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
vjfBAXd5sWmC6+WsVEPg0tlPyoUMdrhyv/eOH2ArqqIuOX7HsCybk0gHRonvAnWu
jdpxVYM/iuxlY9+HNU5mfQhr+RDIdVIGf+LngoWYwn2mQKIvSWhjtQMIxCL7/WOq
h7JdWQ/1SbKAn0yxuEb+OeTBrZqAdTea4k3Cr75Os9vD/GjlG/ndqc3JVMFF/LX6
7lMZA7SVZBd6D8hBIZxN3Ku6mCdyFUMP4+fqWz+GO9OUJNiDu2/wF1RSDn7xYq1V
13KO+wQzNphZtKM7K6ukGiRhmOn7941ROkg4200n1j/gN6Tc7tykxha0rDJ5KwsT
aW/SrsPyhC1M/H/pMDKFL+RNoVA4ddBn6Vhu0zTQ7P7YpLXLudNiZWOhn6tUs/aO
xD1uTwP2AfcP452vnIxcfhphbLebjnQVZwHi8YopvrzY7Taq/JrzbyNQOE5+tsEB
pV3qslr5D+1iT86rVjp1NXiAXT1S9u4XxA6s6etKpgXTN0JbRH6vFRCQgZo05fwN
rAqmarMxn+eGiyaMnmO25SyXyCL4rZMqt+gY59LEPyDuneh317+msKVroGPjCMbh
uNCfSrdbJnL8V2My+KJCVhX9uDqG3NN/LZgtvFCqbMr/3tCNbtma+VI6qNuESkRN
PaHqbbLB6jTyhqv3Yzj9Ii48cs+QJMeJROnghpqeZWdw1tfc4bB98SiGMagMyaBs
In36/x0EAqk7uMoc7earffF9Q8yri4yY7af/Gy5EZCyJ6oKsZrt3sBvuw/9fozCS
e6UxQ3J2tT1Zj0KWHi3Aoi/mxSdtwbrUT3qMdcETlmjZF9CzkamjGGMQJLrX9wpP
Msy2EM0RGnnWi9Szw5CCmOMNpL7zodtADcikirHfXlCSGlLRjQ+SSzbOyJR6KsUy
kUtqF4LYCynkX6VjloQL97s8Me5Ngt0WkPceJDSGvX3WxZam6Bu+c2n4KsCz4JdL
7sz/2xLjq7qMCGyXqtpGgyR8rze9M7qzJ42wlgqLRfnpOHb4ATpjR+MBCwxKO0j+
C2sLDHY8bna8T+ls6TKWwgmmxEoHb+P5TyrkQLylsfvAOoJ+YzAXyxhP9BM7MYv1
P1nok1wVY43U3NoxGeDSqcAcDyuaBufG/yFe5tlrWOin2Fg4/m3krgqKUPk1vmfn
mPl3nuDcQbcPWqKh6nn9qO9ynsvRBffbqM6oxCINNnTjSUVD6IyyjPC3fVl3l+42
UDc2ZjD83SbSIgpuPbR3PI66p0c/ySH979wMIRxB6h2hWRrE5QUiG4J/OrFjvcbV
BIMZx5WJaiEuBaw584zP8JaykdhF23nrpn29yq06gMWgf7BbmwvbdkRR49bTH/RW
wCx/aUyFv4N2IeCNs68N7dmnhmbWP8X3dWisWyKsLXiwlwCNCnCzHFfwBWdiJxj9
IR8xArzrNr5+9jO8AcOlB2aeCWUBVNd5ECbSw/g+0hoTUP71YOcuy6877NrscI2o
FDL8P8Q54yG1Bk6mArsT/ZfJVbQIyAdQ73BJqziuPZLr+n1kholQbYh/MLrMRBgm
jkd53Wf8EbK4tGfcPN7ZlvhzpWRpQBOtEgcoyxK7VuWJQXCaATUiyhgjHotn4X4r
B7VFi4l88KaruUvKD58bAWDY7FdihKqZjTvS3UaKSjXWimZHq0hF9gMZh9kOtUCH
4XvK788kD0Sank/bsWTPPlEx2iQDEi400SUk1l6WIZFb1bbvxVkNT8wUhZcVfsg1
buNW3NBNqbEeR6Pdu4w5WfjJb6Joc380hGo2nSjpX5W6Er9RYNgT2vEYt7xcv78c
u7QTWOrlcDwaq/8KBT2Z2zOd6MJnreOWhAKPRueeS7VzBk9clPw2xmMJ9pL4iK/X
BQcl0Eu0C51K3WIAFiapb2TmU5y3XHI3/udenuvDY7U031ZVa4bmdLdZluaOExs2
jYfJEgaYveGuzV69bME3djpapheDo332lq8QdAAVckTJ9RZ0VHLTkwQ9G6eJ1dya
dGMJPV4WUaAPJ8H2hIPYGPRVgLx1CRTRgw8u6j1Cq/m/r5RBh2beLZ8mjchSqoCZ
GWSx4m9eoRpb8JyqQRTvwoah+AHlsy3TpGqg2Ep2QjMtFRboZo1rjTXWsR6GZElh
zbZR+dguzL0RomnXtMwKJj8LXLWQTAy/l5QyculMP9SXLPWP6QFUB+U6U+GFpbav
PWQL5tLeBRXJKyIJ4msRVbLFXIDsv16VwF6aLiFxpCaWrHYxLWv8RD5krJwP5vmo
PxnmYVENamnPBfR+7hcYcYoA/bB2miM51vUHlQsmqPltderokMWVCKNQxNiyQtQ2
vhQDG0pqpDO6/iJTqb4Qs8vr3DiQyFwIhx8LqQbflyzhGHGP8cjhc6LzmQ+EI2jT
M850rDG3YhX/hhF5vmMwdMWJGyujLn4QCKhQQO+gfdD+hE1p4dZgsHr1SMt7ZXw7
rU1glzuHt0x7k00lahANO73WTfz/x+uiqw0fjUyMmBGhZrEIyBnWCKmPnUtcHQQp
20FJKsIJ5Ay9DPwhzz5kLKy8exAY91SZ7TPDjpUplvrJDs4kVkkHSKomY/jEcnYu
sJmtGcKjIY3O2m2mo8Qx1WxdTBz0XskISM6QsQ0bmd0dTlnVemn84fPKPp2VK3FJ
oFRH6QLPwE/prIU9WLFMlNVChWrhO97HCd3alUIxlgKdOnC/fU6o/jw/HWm12ARV
6dC71lc2dRoWvCDnnPZv902XHAH6EildgdogZ+LNMPOcomFdILKh+3xWgPTJ25+n
Y0jMRaad9xc65KbqHHoWu/tGX4a1rWAmj6KRJLSvlkilxEfSxOu2UJ54yf0V4I4W
33IuPn95RRbxwvZ8H/GaaE0JqRthSXw301khN0V99RXrgSLrf7xusmEC8/D/d2Ab
AYx66T39TsuNxZgffD6Er3ur2Lw9loz6BEa+skeGdjdaoiKGi/llXRiEsBF1KiK8
wP3yrG3wV5oIzA/TT2oIAFvESwNTMDC6iPPfb+w8npAqm8VXdzyoj8nA0inyDa+q
TAq4rKcegd5m4Bs5FSLXNNk0FaQIPkgBh3QaGLIz6hgKAmJe3uqoS3U0hUxy6+pC
nWOFLRldvk0A5WyWfHuKtqFqmdnerM2WdwjWnpfgmfu+1SyFXna7yFS8KwStxvSU
Rf0YljbeAQADyxWg8A0UurgASSyDPeDx3T5hJBbVqr5iHvi8hZ9NllKQtYtr7cHR
BQnGCYhA9jNlxM3Rl80mEo+3bOtxCnIH86TUWzfIxoivaz2IC8b8US9T7O6N6jiQ
DGHZ1iGThsMWZXV8vH0i+eHNlkcQsuInIxPc25rTi3PF6sGnFi5jsQMlaEuE+he3
a6ZKb8Bdi8TUZWpDu6wmcI4j7eRDg6afEXcTBHaUNbB/Zhytls7sYKFQlTebV0NL
neU/dcMmwy4NKp3K+/+1t2ksu3EeIJutVzIozNmi6Tn5hWlWnAyX32nUxuk5+3Xb
cATQJlohjTr0SGij6MGAzuKDZsXGNFAp3UBh67Q7lL0gqXhfcS2I2m37ouwayoHa
HA6CVU/ytrX52YPG6JnqJFKDUWCNkq6AIev4YTQpxDNHopr/mxPp+4TMvnllCinP
b2NHxZZMUf71aDjOIiLPu/1FA6DS5PQhfvxxKIuQEpFCZnQMSvf+evRxznGaznQ8
u69FdY/ikckVZv6dlW+x+PHgHHonhlRhU0e1MH4y5kiU8wXtLjMHgKpQQIcKD1a8
rx8QXHcp1/LdsgoUJfPSUeNsssUQK4QvgWcegA7bkRiFV4q8GGhewzjCa6H6AUwD
rmA0SQ+4MozaNB0L3F04YmOpvwf9vQ9AzYGUWIwDJaRx8ZWHKN73WBBA6nyJP8rL
3yMGALM64+bYHjLF8qhQHY7rXIQTTyEmg4Qj8fcxqT5VmivGT3a9J1DOCUgfKiZc
JmklIV7M88FSsq4fbEu+R6Ev/Ou2Xa3UsbeKJAlrCngq9j0IJNhQLeNBJHuzYamD
CjbkPmUeirthuV1qh+jeCvccXtwCP8IBF4FkmIJMjPrI+u0m9HsM/6wMwDHyHeEq
fy+uKSvO4x+ddZKz/ANEkqHEXbx1nAMlpnD4vT4TmbxNBDmpvgkFgCVBuqq9TUBt
2jUjkZ9i6Pf3rmKQBtHoPfTXEhSlT79IwD6JZsGJjsaU3nIgk02Jyu5T+qkr4oiL
3veXvbzFU/3ScuGeawWIzXteQOFiFJQSkDE4xX+5kTx1z3wNlflx6Ys2/oJDe8Tm
8GMaRcfMJsbgXteqqKPaZN18wizvVZ01EtMujqPB7glPYdcpgRL/PNTSyeDlqqjm
K0JdZS4G/rtqJ0Y/axWdoEe6eoif7+HtJpHySSYO3ssSMF2cLvc6Gl16LLU5tMEy
fqtUYIxWQU5J2EXBllk/XF9EjewZ/eFNIJvBU6mrl8c4miVaTohhaHpCojAFCKl4
IcJMwyX/EpmhXy1nhOsa+Ps4V8OtN7WyFUtiQAS8NjTwMqM3XdpIUWRGQ5sIt/8e
nn8xc5wAT0n8LyzCfP+uXhRZpjIehVKhlgvTaPR0Il3qO9eSx7LtbkckCoxOtXck
ihGmn5lv6EAVG3q0XkOaoQA6wEmxnTi8eGEWZ3FyIKFa4ni2Tadm4uPkN14a0+gn
uBrHtq89VGh2IpRfkyAHVQPXaNvQWq6Qh1oE1bPc5HAq4+dQpwb4h2WI37MM6sFg
kx8spWuatt/S5/TbGwmgrmf/KyKBnSUbMxWz+FfVDkRHl8VKRh3lJd0LQ9bDqhwe
nymdxDe40qfI8tIHIHc38efGkDzTCRu5SH2nwDzMehmJc+GAeIt9C9IJv7MF7r7C
PnjD+A4LUwWEk7pyz9kmcPD6kTWW/fc+ZBoraVdVPsYV6ygkT3gp55dlywXJOp0w
xOGmjMiXmSZ8kmSClXCipxKcQn0rW1WXqsvbtEm6F+icj+pUtwyY0NfzynUlfWaf
yrPd6L7g01kGKtOSZ3jOORamDU260KnH1y5xbMi5pOuIreQ98cLxQ6xgThY4evED
2XuUK8xJeuvliUxtPmBWBYR0hxuWe2lj0XepQswxAcoIsAi1MCJkXwD/jWTFEuYT
KtK1gAinqzYo2hHHEGmi+hJ/tOSic6uc8klbD3Epz9PCrcXcSKAQE3V24sgzPs1C
isnX+n6Sn2M2pTxIW+891XHjo7eN6GTj5ZNdiVWZPakuIXcJ7bQV8cH8+S8LUY3Y
6k1qDwo1ojwc52Ql5zRAVhJGTAmOOj0cIrYnxer6XjE98fJ4N3jqfU2fkj3cWmY+
+W7XzcjJQMcLBP963U6smlZJvORRNJ+MHWmxj8+YHADvy64PpBAviKIggmk6iVV2
mbxTXUJYFxST+jVd3uNeeSpejJL1MMj7WTlt07rfYfey5z6VZQTZ1J85yn4KzBl/
j+mFpHHWRELdUx+38P6S7Hh/SkkUKwGm33PnncFccViliDa0AJ2R1ZbqDEkC+7lc
T5o6/rYYfOqjtqjtnCtd6SCrmii3N5v1wYEGU4gW2jiJ9+Tdd/TLOH2vMUi2pWX4
JYx4tw2qoC+/LSSGyxirUTP4zoE+Wm1jrTNMRa+vyyNbf5QBQO18OrAnfc0GmnE0
NHBrbGGEkzVsZ0hR4K0YkvyR5Q38wT4f78vVj36bOtzPQIEq1eHmvKGUUPiRYIsj
oY2TUcWsSUUUxtPvaLbryNJajw+PIPvd7TXysFCoVGI2Q3i3G18HZ2KVMVInHQ3x
nXAorivaIqAFKz0SeBZXMwxt8GsGt/MEfhyjgHJly88lAkJAFUD9eYNzFbXtNw1P
cQVYVulqC9IvRiZLsqNhuv8bARJI+wkAhKoNY0PlVtT9C0oGgCO5ttbel5Q05aQK
evVigZLPTa9m/OmP3tSapMBVYe0sXpYb7ZwpOxB7eywvM9BS57da/q9fctPKCyRb
/J4/QhbUE2e4EpBoVTJygJu0VW4kTM4WvN2eXhIkvrucpi7MPb1WG4YgVqkYhRE+
gSGPS6FOk8n878xMbT/+jiGoOGgzE44R7LAm+LBnf/khaIrPCHtgtNkM0RVeIbJy
jLbdH1a0/6j52AGo3CDbmusq+fR+y4PofrxgtvZlkXLLstxqCOnbDamuJhJwSfV1
baw/Hi3MG7eSfZGVVGZW/Zx+PvbXOZlDhrsJJ3eIDDJzTeeH6AovffTj9OFAgPHw
14bwo0HO0WIElqYA1m8+QIQDK1sOjGrDgIyf2V9Pb1XJqMxExW46gxj8eDHpm4Xm
8tuUFnSd+FMpf4PzRajlVR0t8lonzStOISiL/cm5LKoDeU7SPmOPT1MMAWGVwVtt
nhNjnwG5Z1H5Qpl/rCJhxf1364dBB8Xey5jrB43Z19xM1/7CR3YPYdlGYm1/MGx5
F5jEaN8oIqAWAoDRyeFHgHIe1y3gHmQSANbCLWJm8gnMSyRUMWXu9iniCGvnluI7
Zl2nwnJacA0ywF1A2qsmjlViXe5AjilhGCGdoMZITuIyG6UyJ5tKkJ1WzDs9TSt0
uuBkV1ihe76tuqI6J6uRP2KKHtsCEQdsQj2s/J4B9tBnbvZxW97YXD2ZLSJmaZcK
KBeOvwycmDdtZdK/gxHZtsy08R9Vd15dK6kjhfNeE2DyVvEoE1bwWUP6YVWg03LM
BNoOfXxYEUbh/WBGwIfDK9wZaHELKAtA76V9Ut49sn2kKMecI3zCI5HUJe4Hf0l/
33jpvk03cBvPQ6bZuGJmDxLp2v39azCtg1/OEOO1vCabWGbKpBkEB2AdEHVNoxLG
J4/Iu5XAazb/CXnLJZaIAh7WA1vNfDw96CiAcvp+XxNYVmdFjKivrDeHAec58tcz
U389EWXjzf9EvvJIhLvLKatPXfyZxv2X7wTV3bekfJnITqyvJfgeu1ZB6kjLMW6V
Ef4HYHVMtQHOCCBhF4LL/qTjZ+baHwM+z0IHqXkOcRqIzTurRdWSo3070PPqod8q
D7IIzkAECWRoMqtGD+i3FlOTbS8+c+Yp2ecj15ZfOOmFedAGAHsRwDveY3QZcKht
tN7q4pKJ1k6ujNYivas10Fcc9L7417vh1e+z3IItz3qeGR2X5LEBGh+5VGf+zcuc
RCyg0OxX/SoJMGLRNAUJAhYiwV7iAKBkCR03V6MFR49hIZY0sBlTbZIP06iNzwtt
uQMOVv/+GsrYrjTogyoKDNghgICNbY+jExdJwt9rNtFBF4tWgYBFmIc+Avo6tOxN
uJoYnl1Fny6/cgARG6DJsTngsOk+ShSls736L5INLjiEjPtoB90rizdzlO8e9tyZ
65qBhtOrXBM/2n4iNXm2/01UOnDWZa6O2ZjyvFKxBvRJOzXcnrnz6cHUnMWdxyda
B6hqRy8E1dUBcqsM86S1efu2WWWMANaYqMP/hMUbA+d9fe8jKKtrLWBwP+ipA+4z
codMyOcaWcGxrJnn3wJ8J7g1k8D56zkfL/f5cOGqNtVEP8N1BF9XZ/Yk7B70rub+
WKNjMwEDdj3jWCBK3sWA5voWa5+GnHjxDqZ8f8w+nNISBIixOK/sDKhL76ypy1dT
mdIW1PpzcA9ABfa0UhB/14DfSHcfUrqo2Y/x6aUWYG4sTSkuSqYCTim+oKk6rUU0
rPB0I+Bap/WsebdVblJscnNRf4oIYK+lnZZ4hLrPZxRBr3RlzI7FdZjo16N1ulLj
LGkexNCjEHegfDUiLSXpYHBpIbBRpgkFbIoGQrrb2KdRjd7BEAGwlDzv+mJRuMpF
9HngIBXTx3ZtGrNz/cQ7ocoo0NldQ5HKpXpVzcMaDBIZZ0auC8MS4HLyGid411CW
dOQiJGje26CtCzULEoDIEMRVTo+O60uWdeXKLnOMNJqqAOLFXw/4EoVcUGlFgh1k
b0p1k2URoaKsz4oFczhtbn1Lj0BxoZay6PbZDpmJ5/1C4K6SiNaBur21K0XnO8fC
hP+/I+dFk1/X0NbpYx7xHYRwGq/+rEcaZji52Pv0l4CvRQ9ikwuUl+E0kABYsjTT
YA8WhbFctJ0MKXUaX4s75dLh1EX26Jin7cvqvaKJn3k6eewkxwK7V+7POxgYczbI
t91754KjAQlA+aQg4VgC7ljlCJTN0GMkVRQl2BEr2FoYxb8LG1v/Nkp5PGtme9Go
O022UXlLj/jJ5zmhjkbCodLyf3LulUUiQKGgp9OZ3EtRCzywMS0s0xs8Vyu9V19q
kYlZaegQ7y0GHQc3Ig0ZN4QtriAudqBwzx93PkGYy0MlAipEh37cLDIAWKM/CLwo
3cILpBFLsz6I7PZm79rKj/dCuK/k8+VrDSwFohxgCmS8wD9Bkv/8mn0j81eCQoAw
d4WyQEMaemCsTeJ7NTCzA1Er0UGMdZq8tbcOnUChvV6o0HUjUJ3VWrRjzaMTdoTE
Z9rYIcaGeelKS5/Z+HGZf2oTFaOTfFAWCasRnClOSRxs76x4QKGZtr5y2V6MDTii
bbnAKfXJfqx3QN7X4RMZutBSXfF7IA6XyIJcgaezE80v3xMPm8weT44kw5ejh7ND
pGysYBhnPiRcOfYw4LDqSn1TnDXQKJ9zkd51B0/BywetEvzJnCwaq7e2bZMae9Rx
54m5M9P0Nl3cThwtiN33POAoJlDEdwgmezSmL5z5oWwKjIlMwY4BGxjNRmOzJcVL
FDnw+xOapNCigli9yyg+ahRH8cuEXgB0cSCUTuGva8112w/+LXotygsKnUxp+BOI
4gwToaD6kd3MMUW3crAH0SncxLnMP3X9hI5/N9Yt/j3tgpCV1HRcnMbgHIUfFQT2
OK8tkuCBCb10WwTQMY6xkwK4n1tp2Zb9vEMTBiBjQMZHa86N4tmKTJY27W0YfdJc
z8P7Y2r2jvuOx/n5mFAb/fC7Ab8f4/mgjE/p8Z1EWG9XzgjJt9esvYCTGH1+cY4V
IJZAijAe0Vly0axiDS54lRAA4NLq1x3XRQUObiCPt1R6CiLL9Ump+QeWqqAgfCNq
hh+4Ij4pTIzijTeBhv2ZPmASsTEnpEjlIp2rn2tfRzjHIWbEmiyBXXeo+6ItbHQG
vJvC2tYBhy+R79Yzumj3H8pfrlP4Lo84K5eS+DE4hfgRFj5g1xLkBpn32W3dajyQ
3heeQxGLkLrTguNWbZmr827Ki8mTH4aiOzu2vc5u2FhtUiuaTaNfpy+75CvjK+LV
1B2tAqCWv9H+MuksVePqeXxEnTXm0+tXuzau3R3lkG7hkz5zKnH0+xinYNO166VX
upsoxMbkEELGDBv+D8tvZkdLROPKdian3NYUjhaF8U4CmJ8Wjb2Hz8qRGEdIWw0J
nghNKxgbJ+/MrSPlhpbLO6k8KXUsyP+MbWtmLNXal3XrzENtxl1N5YJFWXVaA0SO
JYlgnKpA70k9lqVA22llYJhsGJYM/h8qsjgkjuLZYVESr4oYnHRiDrOL4Er1QqTy
zB6gXSEnwIv6JGamTW4oZ0kEH71XMlAtG/iHsMpPAVB4F9DOUxHwUHy7UXdfcgZ5
yxhKSqs6G5wlykW47SWKV77SVbNPpQQR1RcEzvkB9iURYgrsMkVq4QC6kcg5jjBD
hSy2PPmG/X5QkWG6PDNl1Jd6jeFZiBdOjwWsMM6AjvsHpTtD6p2CTNrEolAfIY0w
irKltkbKQqYnbov89M2ixBN29XaeY7HA7UEejWnAG/1Ud8DGtQ40tSXb60IUxjf0
LFOtDp+1HQCY4fkCBfk5fC5WrEsjaAf2UcvU7Gi7C+kngnKRRKV/86bnAdG8wcul
n0FUN46tZy+luwm5WFJFmnp28AE1QMMXdVLfz76pJDYtF0E+r9fywDLI3fLxFJOg
9aYAaT9PbT+ggDGF4+WO3wiEWGLS9NyPvImZB4LenlOC2LBJeZKantInCIqT63Gi
FAJs+I5V+Rlal4xaypplUCLKvthD+xbIueW6u5TxAUJJ646TYpoMmY7gzLaQu+Sx
tdV6sNaRwlTjBfsFw+XB1VlynejjU67JsbHC9dorklLZXf/KuW2fnsQvbtLHkP39
WbM2Ze9CwUMMPpS6KA+FlwfIqUpvxReSMo9nNHIroHITz4Rfp+Sa31LRLcM8GDfj
qG9qJa0bGPZ2jSWMiePMaUYEVKwoZ1AoxofH8zD4U+6qsDtwL2AYhEYF2SedsB7L
kE5orUbaT9mV8hBDGSrLUjkXb0RaVPEwhCbwW5f4IggICRJIINo6+Gnei7XJes5a
Ai17V9tUMSY0LFxWUeLSSQ/3IGs/cvY6xAmQwW9lvOqcZpnKFAecrIL7F/6pBLas
XsG7h3QfxsgiEobHxieoea0QvOOgaMox155V7w21V53Tv2D2q+oWVuiJ1mv0w8B9
br+HKMVZNIj40KqRMc42YBXD2aXqRZEinQwFCjK+gFx5SZKENQskrNI8OWL6e1u0
AxrQRq9KfqBW3Sl7c+9NyqkJ1mCGHOqwqioZmITidlPdJ9gpnK0dRK71HtCDWomY
6PQL1IkItKAG2fVL5ZF4mDC+bnx+rbMso+/OaRqRnNQkTm9RBDulAay6AZmNgF6k
2yAZ5E9wd5AHKik0NLvTzWez3UpdWmxrlAoVoFr7gLUjkgJ6EH3jDISZ0jCBFwDE
QrvtFBCu+iHsLdGRq+3YCaTH8eq8mhhpPVd2yLfwfr0I6rswu2B3U7KFlmnKaAJx
xZhdHB/mwsIs5C1xi2XTiXTi0wcznVoNnpnj+JiQHQVw4Bb1BU0yVHUZ0DdRxHZT
4ElHBDbTbjDRyALft42VfHFTtDsuOgZHtSQm/obaFowZunHsop407CJaIS/7j1zX
pZ/GfTwQibjd8k1CkwEpQqELLvBAYtLU6VoeLUiwSe1zi+h199sjN3SKa8lYfj/I
cy8b9UyaNrq8ZosLj1Wt31Hwq9bL/5m4aSWLjGHAGpz2UcpoVZW2OsZ2UBdZfphn
GYOOxZDhx59fB0lO1XtVKT73B/Cf+SR2Gnniixuai3ZEmuBRvt3fDsXz9BpSBFIo
yfUC23ZDsvU6plz7maTC3SFk64rSyY9NNCDWRfY2qL/PeudcSXOzyKFiSGC8vift
aATgwqbiUQaJc40hkECYLS422gRZBPz2NVi7C4Kro/HNqciMfxgECbY3eLkVdSYz
pOtq0ERL9uTVV3K3yCtjeeQWS0M01qK4l4r3Nu1k8GqWexZ7iPkz6201Rj8c6OPU
kOusxrlp1S3OMDDwY1rVjLS+G1fc+O7RJ+1gm6A2MDm9ZXZrToqhvuqr7PlXBHkk
Dg7mbJGo/NQmz4OGHSiPOrXMrIlSg1rjwcSV6Nt0pbr0GPh6dwPQGDykKi964rwP
mBNPhFOl1b22VIgPjHRqExZkoC2ub8M6iV/ogczWW5c2+EzUYTbLcQUJH+oCUUDw
HZqBH+bGyOvdg/icOdmeeFEI5sQhqMutmQh3LeqldyHE327VY01k1RV17VSD8rcN
4HKFJ1LlqFQhdUPkv3W1BV2qSnjqyBaw/JTFob7RmIfeclNYb2rVsvAEYPquOUUG
WtWdDl1Iw3/VekQEM6h4pPwG63ZBh0h1gMnhYVvnzNb+9Uq4iFeU7817axjg+WPb
twmdsAZCR9SuwxtqwGtEiCQ5ShOrETfgM1nwSddkA61T3XOh/mGY4k2dnq2H+ZWJ
RyGFU7nWuGxKfL5zCA13tFSxff+L/Sevd3pwMwWewNoLdJfPDQDouT9qOZFvoFip
yxcMUvG0XwViBrtpPNQL7TNlWE/N8MAHynvu/SWaJSOUHgJn9kZksGIJUBSErfoG
Tlk0mEHSZI1WNP+VLzcC+Jp65CQd7+kC1ei2PmqoH8zb/zO/demnF3y/AiXhzjHP
RsUgMb3yC+tYX3M3C106RuKzyfoT7LI/U5aFzbGwhI2iVTztaXlwdaqDGqRsfItU
kctnoq5bSOMXP3s0hAoUGHQrC+QCViZ5uN3LU9Z1A8yuvMEv2tmVOXvmAgWodFZS
syL9uK44KBeYR5pa3IQdgIi/jAEd3PEiJVF/bobG9SWrCg0q/ADGaP2CNs4rz1kN
cvMsmZhsmaQPUcBywGzrhpWCLXPBff51s/7sWV9GA+3OUjqEXxRnbNKCh5HGrb6A
j+gdzoNphUV+jpTYulvvv2NsGJOvw/z65obvk0oROl+NABJUlHHm5whdU/lN4l2U
YbG7ctkJj/aI/EpEdfnk1GkQcliXWWkW7Z1g9kLF2laf5o0oWF5vmgNAqTDG9Shr
aOna0yAGYvMHVw9q7SLkAYDLhWC6D4G8rJ/ib95DojqIakvkaJNTgiX2+I+kI7bV
ILbx9leKJ9qzGEBG+B+kIytX3l8l9cCO0PsQKFqMDPLhBTTol5KY3QkODnYEnhBm
O1g55YJf/5/vbjtwE7xnB1Eovhpmz17c/KwOenYE9x3CHOiJuvnxaMPqbhYMMUQC
zr16cghxWmkclfMweWWhMiFJBMSm2Y4/BCDVtzxHxcfJUZzz0M+P1EY/9CQh1qON
FPc9GkaU2r4BZ23RaYzc+i6x/0smWmlvtWyNrlxXyxpYYCMwQNzifUTvZcl1S1Qh
P7XPh9Fu9+d3RV7BLv6RWC6unK8OAAppsGUnHt1OfpU7kSWXRXecjk9uQDgyyxYP
JAuXbKRHshjwDks6Cay39oZ3D+ZKC3Vru/DWJHraD9SmKfEII1zDtncXeZpRfb8D
AWh/sSD4eg/J9LxTAWq4jqYFh7WiSn6LIhyhL3s/Jt5JzLHfAF/cF8TfhGBZc7Lk
o6CPEWs5sFFehQOdFLQOj+JtUW2ZbPrd3bTDrMsPfYxRwY1O5tWgPX9a0/28cGqp
Uf5TlHMa2GqrMNYHTWXVqjaORRdGebDVu4IBenWgRIJq7rHIENLHg9iz1e3jVtZA
bbHOyf8og6EU0/Jd2qWoWCPT1Gzf2doOxnHXwZqglQo2d0fNtboNmH43Eq+oa85D
P7xPWMMMfNusgtCZLO9qF7gfArv9GPV7JmuDUlKwMXGjuVnNNbX7NhciiOxufury
VwOdCYzIW+U0EpWVcf0VCOSR5K/avrSJFGWxPflk2Y+mGAgt2N4kaYPaqlsDigfW
km79smNfo7gjibhMj3wIdIjhNgI7fMEEhBS6+st615ReoqtWSJGPWFBQ+b3s2NTT
3uFiiwT3Gj/zKEbeB7GRfIa1stIIGBjVS/6yqlgkBSF+CYt+sK4ZqtqJW2hkhREm
jo3WEyUpfq8fh/tKPas8OVp7cQJya6hR84cNydKkjN9uOyS5hTwNYSCZf1t192E2
kmyrZ2xAYOb07w3vSN4zPWXAXCN9KCBpn8474p+w1eReTs0yW9a+yeVdTLhUoY5I
kiSWyXDtnnLbcvxImaRLuTPnb+M02+NEsEnfQrA1mD1uZpn2Dk9s0l7A6yftS1yG
B/U6j+T12G+2p2FlF5CQ8ON8WPQgyiofEwEfONH7ZorDoquISWVfmjCtEOG5nLmK
rdFPVBgW5+A2M1Utjx6UnVmtjBh6yOYqpHgm9dzm6QTgi+jV2l2YvfPJQZyIuY4W
Y46og2Q/T1Hjyb7rvzQXK4BJa2XRPCwfegkCwvSyy3W2yrdHImfmaeH2oGPq2Imy
2k1SmbRZV+NySwPs8/tJpW7VLia3GJo2XGDvq5A7uBflHOe7FWZUfEVe0hVKM+z9
vCL9R4IVJbYCZ91My6gfr6ig3MvjrnInJd+jKORd2MXDm63Stv5rwOlmE0tyA1Cs
j9cnRT0AGczLJ8cT4rPbyD+To0zgwTs/lyk90/z4vecQE2aCEfE1BTpM/8rnr4on
jpZzPiINJBUA7wMODU75nBFw9zi0DPdD6YbAaSxELWrZl0TJUndiT24VVwPlrKhw
/wSLrJYbtAGmRd7KtCFyA8M7tW3C2v0wC87bSu+Tqx+TS5KYosTBimZnXZ9wA1JM
Q38grRIOj7QcyWE62zjNFtv3PG26KMbrioVHf8jChV8Fexv8tTu9HaKdkRhGpzdL
MeQBypi2/M820/gbwXfBHdQzo7w50mDtFeFEIohu/UVAikCWWtvhuAema8zHfoZ6
MjuRVgORVeVAD9/ImfXKcFwNnM0tfbWHMYkN5lVEpjJ7I3cmSWue97hPhIIjXldl
guuNfY2Owo9fyHpUEurfmiTXoJHCtWKlfPEXjwSY5p7RJyLLJFepo69a9/fenYUG
AayS41nHZtYFBbqG0yoA8ids6p7ECz2lEYZ9sseHbMxsXE/F8cEPlZCA3TC/Dnva
kauamG+5VUxTFGkeJTNJt+1tnEA2M7OGCXM1RCSY0gnCb6fjCIuLRAPN9YV5tuCf
sfUo4nijA8cFOQgt3kfuphuhsSMAUjRqnu7YqftXSXiAoL9QutW+hF7Ww/BQA7IX
SsYo3/mQjGq4UUag5kjF/O+sG7xE1tduVCzFf9XdvhRKwVq0ykrAyzkf9v2AZv3/
sO69FTR4f+RTP28GUDN8oKUFE2Q5HBlxj1kg88KevEuAKbSnrdzyK38BJEv+d9TD
t5AhB9coDPuqsTUq0OSNXpPpXIOs8b81VlyHROmVGDDyK+pkadmvUxRw2vs2BOYY
iSuSXyY1mlqw7qKfPhaZLIp1OtRljGHsJPyZecLf1r2ojgLBNNCz9RA/zKr5/RS6
5+1SX9exKQrhzkJ2pE8V4S1ioBDQHfBHx0BEvlpcS6Rv40teoVuBlyC04MxT5Fzb
HSPwhK4IlTv1/mM2CEQvVFQKGfuGL6YJcqLzYMDsTWclnFFrgYglajCl1elAYZ5j
iiZ+38vAQiTEgq/BvNG7irGTsFI8pU3gHlpldCmIAYLRnq6oHJRm7YRtE76+J21W
69MtQ2DgglxFCMyo4KoNFt/yA6hMqnDtaz4sXR+0lGmVP0JOtDfAtwk+gDcYp5Ab
ef0w6hQxGeYMPv+T6ora6WmBTcGwUZhnemdmPgaXGtJ2oM3XnoR/iZNuhfRZKGSw
4QZ7cYR/VICdXzzmNhsBMyLe7djiFmatesb+pQzbsO7l9A/h0/5cB8KP6ceqwJ+a
VoHPuQh0puGZ/FKp4FJGa/Vov9BT8z36xLSwvLdQ9yZlfic5leMsTmypy/zb+YKt
Vu3kit4fdUkfjoR/Fccd0gHUMOvldvEP9ccrqxSBPT4bzBQU5oundT1emBl0evqd
YWRMjbgkMzE0+kWO2orWgQy0kOQFTnBtfoNJB4jkOYNSCHzMwPIvEpn3AfOGN2XK
b8+RTZxUvkEcw1VInyZeBA0WIxX1XKacDO/DBMR+rtiTymcT8DJSqUWRlZUxAqo3
9ESpdD7Nr3i/C7YNbNZsv3qmc0y957b0qfvuMX+DXpcHuFeYNwcVZyRbt6fxPvnZ
Zue4TAwkBvgnS3aW8h2cIMMVB8zXawiuTbjHIeX0+ZhQ4KtFn6fRduRhZANaWSrk
d4CMJEKvLui7YdlXEf7EGpal/4azwDBuUifMGHB7Sx4Ti6p4dvuVN2ng215ZpdMI
hvYEfX417bgR98aTCKZEiI+K0ugKnqj6BGsAsfva3jKHo0go8A0v/0BWtQx76AIj
JPIqaFRM/jXbaQ3k4qaN9ekV0isba4/F56Obk34acovzasKj0iwc3OtpMTQmr3f/
1y1kgtPjIS0ilesGKlZT7A2yTmOfuo5S7wXiyfKpChmtuF/fNxCGDzM36PdZfcBH
WQutch8DFiYytrKFOeJb5QtT0oMoTz/6Pwk+36uXSEGry1Kee9rVhFaPDPQkXgr7
8OzU3T7TgLrP1dRPmgNz+By9ZFg6HR7JzKguQjmkcZQjppVfRUhKaRDzdBPnSUxX
obYpRtwNQCA1vG7rDMTYAdQ+GWHrv0rWkNMGC5J6cvsJyP9buPCUdHKjVwDIhhEf
jhsZTW+lM1LBtz36l16Es1qRQ+Rq1n8wT9R73kbqvNjfO81M52nKzZo5ZaGW1KOE
O2QQthms6etKePpP6zt2B/TW4R5TZar8M4DPVjLO0SkYVzabtqm9vN/n9rYs/0rJ
jgQ0nCOPpEdhFV+Glj9JdR3ThHa2aMrhhrYDkxP6vPKQF8iK4FnRidf2sX90T5XB
TCJzMSIU7770Zd+YTNvoYfhmIpIsjK/wBwAHUXsOO14AqJs7Zb2HvF2gSEfQbe4u
17icJkpvuUOOzi/ngQH1PZkoeXWwe+laITc3xVQvgUjF6lS97ZHqPwhTAaUX6xuM
vPFGqrk6CBzar9GSmLl0DZV0kl5qUNah2ERImHK9LX7hmeB5/QF2Bzt30PrFxLme
AUOIBBOMyh0UxAj3txt3vGYWenswhybn44W6FW4UUNNqSW90SoJRF+qLQrxollQQ
6RF0gDYDC0p/OW+Slzg1mzW/KMJag41yYMNr7+oJGWm/AK5St7g3wHj3OqQZYQw9
JtJUf3tcq72EmacI5bJU9n2ZZqr08ajcALm//RPNrBKARXy+8aOlA9jpfwrShEvW
KiW+1k9R1/yCWk+ZEHKXFdvQ9uzeYnfuypSdEJAGAuG2zkZZI0VProBjRktOIz9u
4+nwmQoeBaMqZQgKvFnUvxmdMgYFjRnYfSHw9911ce4jD2Tpgf/Px/rpHqenSZ/q
EgYtQg40JqFpBEj+K/x8Ue8d7Y03CH9uae6fl2IoMFmmXlqNipBJM3msgOQYN6CY
jM+fPDX+peeM0Ceik6CQJ+1+QhJ+fyzo7CFEXnc9HMLGerzmgy1c86vKG79K5ui6
U9VsgndodTkCYngGgnTthFgwaUBKH9dg7Q+Keqcr7X61liEj6SxyMVRE0jbFdoM0
LeZ8FG0v9HrWAuUQMyYpH5F3mxyl98LyzK7MMg6S4TGpoGybjR43wDIjIdPPKUVw
FN8wg4A+Ez6P0TWbFuoUmigPocvzXXdLDcFR/bMMAreSm/TEQpyZpIdCXDCoioe0
5xjHvWsQ0t9BHL6d+AGFG0iCdgkta6qoAHiFVk/JSMKdcgGRUzOP8ecJPI0KVb1f
Lce407NAaSSVYOR/+VJaVh+a6uTAK8jhT1IkzmIsihc3YWwCRgeezZtJcnOe8sRq
BULV5dtm/NLA2Y7+EMx+JuaPtULkhI66K8cPuqkN+NyCpCeW9+COM+DEq1VlBgty
0aLAFpb1j98qkbY2DrzmiNY8IFU6Jr8AOGFL4Fz66FI03xAj2GTApK2A2l50S90s
3wk4EH0qXZGcWTcBsQSpSqBn/z1PC9AvSGkKeA86gZz6mcwAm7oVm/UyNCmx2VVR
1CBMGoCgixWVR57CYRoezH7PszCEZW9Sl0ZHksJv0wI35i/CVMjWyZB+OU90Os+n
Pcq/gvLrroV8K4T7pNMtgXhkCT/phGLankPSCQC3984dd/FR/hc5krtHem1IhaWk
2Op7lxirP8szla0JOZa5cuXtF5FynSsBi78HiTacg8f4XBFRC2quzYf2svWRIqGF
6ZkqrAPLWtZD4IxqnoF3Cf2tanA7AOdF23+6zp8MpUVKiMcp2OYgnI+s6Y9YI9L2
gm7yZwqC+yiT6w5lAn2rb2vPpHQNaTeKJQQlluMy3QYTF4/F7cIkBwTIJIvvSpne
POCEHZB6YOoZR2ffa9vMrtIYJ5UVfTlxiCwirpCDROfbXr3up2KBwc5FKDK0mQsc
/7Xv6cvdzCZhBP4+g3MV/gCH8DFVyIyS/KSuc/3zRhuRUFRVY4u0wKP/+79HKPWI
4jgIM/alDamsiDQlpMJ8lYeJss0klV71JSDbC+sNyu0TMvzx2z7eswFzhUYUAf+S
DbQfib/nDxDsWxcgCObdQHscIMVwz22H0wZZdPmZxq0OMHKGHSwEK2dJqPsR2wjy
DBdYMEDYnTRAGKrBnjmLJgCdrPkXsLBNxGLHEQDICF13U4h+FT8JmHjLR7kzF0yY
90orvdVspqhyGSX6F7razjiQnjUpNouInvgzsrSJkbsvYgYuXDfQLs8otzo2LYwz
lAy1IRuns58fW4xv/PmJ1IltCImZJwGj+xOtfNAJzn6o2VI7j8R4f35tvEPLvIK0
Z2aPtXHSrpBM80P57Y4dGnok7gawpJyvEzxUhLk/ZHHBWttDQ5Nipnc7boXqBbRA
6BneD/6tbUcgM+tnNQ6dRpMvbW+bPxqW0efCmXtXVL8+UtA4SKP/qcD1Zy6yGeS8
6isr4TLKIwgAy1AyYbharZY64WBsw+g7Gj3rWUz+MY7eojpOIUKOY2NeRk2fqCU7
/9u/i1j+YRqTMzBH3xol+iMCSSZ98c1NjFEO8N0muL2GC4C5DvmlB1K3YG8vNLQ6
wWSJ0vs3XT5jbUMCsAw+AJ3YUrscoe1QqnIQ+dOvPMq1WLfO0eTcLUwWyVt2sqnh
0QavKI+xsMwOkPmzlbx6EnpJCh5pykME7MurPq4YsSk/Sl0fmkFWdCcNcOrwMVF0
ZFXG8c8upZhrm3Xv+tpavaYJ3zYZCWcHu4frY6S2vLq4rV2bjebrZV0HCWmQqZqE
MK8pwf77HJv4zj3DRLQQAWFLOUVGipkCmTwuTSexMJDac+CjhNON3FHjfAZAjnA/
JZNxWu5wyA3jCKa5x0kuGyJkehOfld7go/vUDgQGQq5MXzJBO93PDEUIX2g+qPsb
0BT/9sYAwQm7DDEmrPqawOSmzHzno7BYITMAykDCvLgL0W096sff0mieOImEFE+5
xo8D6JVNAs+TxXwTiUaooVmX0NZ8LrYquBL4C5u6fE9ecnOos+8CSrX5RLLVHael
XjafldmxRcszaVMy62ujy4PghoDS2SlyK1dCWaezvHb5n7vraOXuoS2d+FCyYwUY
fZz5PxDaXVEqhdFLHyY0eJYdBesZfmM7VVPGeit+B+U7Y/xgp8Hev6xHL+89Ltnq
AJp/6hlvrH1bDPhE0qoHiyADauEuqdufD+qc5SwNLmW5ahqBCjJmKYQQ3K8nDoff
m8dHxEUcjbj8HdYAPDQPA7lIKWC1TULKIGythgHJwPZ+LQgFdE0iaedrcx0Txn1i
XqV1Zos837ZJpz8MZBIzMgVZMzi+zj1SAPnS9bTqXXzOjIiTd125ABSRMUgLO08A
oTSMMtoH/SXZNdEVmAsW3jNP4uV5xM0lA8cE+NoPtgrZWT0TWWH4EAejV91T5s7B
GUy9BswVFx/TpGAlUJaZSOq2rxpIP32eJaA/yNyrX45PW5w/kKaTkCtdWz8UqUpG
P6CSL//otFeAus78LtvNnR+pBZeHEHjVKErbLmnGgLrKSmJn7MFPW2u77l4HXwJ8
pei30kYVT6zXabrbzdWVJREdfdcCC4K/Z3E/kxCcgjZOyiUz3MvHPV/45j+G7dL/
r+tRl4icXP8CpFJRwAaeiAdmCqxRP6RgITmzn3WgvOCGj7EDgU30QT2RR7U7fosx
zdlCgddU8rnAK5uI/rqWa5leppIQ2onxSlGssO8iJ3oY60afaL5TItUq/wc38yqU
EP056dCCPXOOSSqvmoNDXey9e14a/L490FaQm0BA9LYb3+lhChE7HD4vUQ+8cJmF
FLdWXIZeW5hH3pXTGQk13Nx9VLBgEPtdB6PdJcQHKRok9ouBU2e1nOAzztWAyqAZ
piuYSTNxiYSekTH22nnKJuO8jD3X9tghZMAAFj034iHQZloDbe2/DG2IK4R0Ep/N
03NFzoIAvcL1GYQnxdkERPU7X6AvrzSKe6J8dfKmNDqLKnpzMCBW/Ebx+s4O9cqn
EfFZKflrw4j5YGbjUCSiXSqGzX8i7q8rG+FELuhrPXM1dMmAydnNpbspC5k5NbW5
3qs1SIhSi7j5gn73G3FFHqhn8vf8Z5FyYpoOJJ53duRLiyZ6qp7amdA7w4vKFHF8
f46q5Fdy8gOtOHYssxVWxbhalU6bxEmvAQ4FGVlwRTVLlTwav9KAAxsroaJ4ucuq
JQZY2mcruZCgZWp/YDCWojpE3B9/x/yG+yZ6eQ2zcv6tdCMVSzzRU4LveCZNg8Tw
5xVyugZSLLlvgocMkIb8DMVkoQ8weLVwdfEteDj7KpPWAcZiB4wtFGtlDmUL1mW5
SsrIuXfSluUhq1qRmL7zrSo8WFmkL/KrjeNOW8Ufdf7sGNvfnt/F8niCjhikQ7TW
hgBaw0Lt08MwqQW2WfUqqOgRchO+nC5MLbAaH3TQrSss5bI4Bx7h0BHgYpt0nwgn
fTO77H2YKuUdT91PEWn3pdGXBES1dr0KQGLVsSxupuRF9bZlNgGRjXAdv5BBsV3m
BcLR2IuKG+0r/cFVMsHUL8jarCcLVlZObWOpyCW7Xpa8a/XaaRj6hcEONWWOwkQd
7grzPUfFvsV55wqBBhzDqqw7CMU4ePUWD9fEppWA0TKsEub5SnmkPFjRwG4/XBN1
OQbcKqKMm6VfJavcXBic81hXEIxPtz2PSTXWFlG1AsojIxgLYBkFbpwrhObIUxj4
+FnrAwDXBGYkv1h2cq0nPrpEbPt/hfcdX5iKLpe/68eBu0FaGHdwzEvLlxXRjq6k
ycMXlqD5tBdI0eJ9H1C2cja0EIpwG57kPNRHOASzs1Grcp1T3+UA8GEYgIZxC+my
TaQa1hYXEmlJQSsZGjHJ79ZDiOtcJ03zDmwo4kOREmKAtAz4/JOGOlaStditHHIE
4BzkuX7mTSDSib2zMiI1qzLDzcONBztm59Rg46+aZd8nvoVdhNy5ar/KxTiiJ8HG
LvYehEe5L3zrCqH0CFtC0pw2BZ1oNWhpFMdVYGmE5B69gZm4yD5HFRMfjkreNYxT
BjEa43xseDYqJxlkvMpVPwkqMlZY6VlTgloQPkOwYmW0tKELSVmCm/WMDdP2bsic
lpwSXYl/klZooPULXC98hjes5igoikdRbO0dgfP0F/PWi3TthL/Tp0ntAzlPjC3L
SPVqUnP/E81eRsDmgp3mXQfa9uxdID42xrSw/qxXiZ74cN55zaIialAOc6qHczLo
ylp+Y4e3MvPwsaB5zeppmis5XHe3Gg1r1puvUPm7WRon+L/50tflWFx4Nbs/cDpj
sZ3OFzNi0k8OxNh4jUYJJjSGjiax7CBssFfdz8U5D1JxPe2iq5GIE+eLrFoNkErZ
9Xaltyges1r34j6lNi+UdhqZn9cYnVvWgYEaTNtUGsJ7wdQCghACs3rsu/vFXati
zdeAnP130077PSGtIvES+qC10B4dh8JyD/r7q3Ztfd1OcDqwFU3nNM+HGr7My8oy
ErGTUll8GgaRre6iA9wWj79NTPpcFBTMt05i7BDy2FD1Oj1K8vEuCm+/pjaht4uO
Y3VhMG1eNVX96DplF+uk4yfipb4BeGG9yd5VQe+JGNEEb1A1XfSntQWNMQY8nLFi
CqS2LlW95srkd5YV7sFndNgv3vj8pBIOJdlVYgmtEl+9OdaBzO10krDmsUcAonXw
q6fjhVRQBsOFsFKm4nnbXtxc9YRIuzQ9e9fCus8UsL4XkFhZRNtN+u6JaWcZEqCp
iGLXDBg7hL9CkRzyilndzm+RQAi8PHqdlJgxNWdFwDr7dnzyONR0wXN9bmRtq3qE
ib4w8LJD8eicw92d+TJoYj4akzN+niRQ0X9T4XslBrklOTjuZ+5gIU7Rz+ulqnmu
7DQgYHkNItFx6jdAghex8SiLoVjCqGB8UPS+8dziJrN1R71HazixgCcBkKQEc5gI
Piuz8wgcK6TsNDolX3OSb7TvRQsTP/gsZ24ziGF9dRQ5jyDdrG4i9daAOhr5gy6A
uhSxYFaq+6y7Q2pCVF2oaztZW7BDPR1fqP+oHdXbgvFl48rIurVrri5LNUEtrMzS
6EQNpD0SJRdOmg5nm26dx7s1Ul3l6FJcUzPWoOuqxjQNuu5mvm2ADpN+UW9N4447
wIcqDN9X60Civ7NdUZrCAKP/O7LZJbNpgNnvwD/TYNsmfLWfnvlvZrAsQ32vwR+9
8vIswwESiZ0FbcU5bs+rZrLzoTEyihhTZ8lUiasXriUIlpo99MXYX9CyzTFLuTbo
/+5+y2rdtXQ0iiUoP6h8K0uqQLIupwqx1nRtVlERivZ3oBoeTgkdnpXTMBiqV8nt
TjVqY/31YMFQwk0NdwmoCEW290OIoD7KUQs8sUKWuaBWL1Zh9+i/gSmbjMama5cK
hfV0+G5E4C3wmwO3ewaOpreD5zyR98b0hCueeXu7PP5ROkyAhKegGw8bLztVlSnc
epyUxoV10AOuafvigSV0bbOcMfTlTRdESmtfvX5N9OZmfSh5Ly0TLR4AyAK1BGxz
Zv3NXHdeJ/iabqbzcj2kYiAYjQ84xHoiZLpIp92L+ecp+F8oyr5DnGb+wB5yOTCG
mPsk/ewLQaKKXyhD/AJQkUMW7cuJXjvSWtksqqhW7tj8TCr4Wl5OkyYBeEuVGB0t
wNbd1M4UoMUrfhsSz0NEkXb4wd8qCyypTcz1c9oIvIPFetUh1SQMN8XUTvDWKsNu
y8dTRgLZfQjmOovx5L0Vr7inTm87qV2BbU8H7JV5gM87SGZC8HarGAXdTnZeoVJZ
ydh5TKZs6LAHdmyb1Mixeo8VhQ+y2bupWvnPtaReaUTz6VkEm+sdvz5zFWKyFFsT
FpZxl4y4C8ojRtKst08jjZ5wDr0NL5beJDIHyaTNLETWx54CEj82ilo+hFsDhsXG
VZDFQIwjnKbELWXI+B6lujl7FHOsPNqqDaJJ53CW6l9Rr7Cwa2I/fmChSQsMpUg+
shuOAaDNLnTH5NeycpHjFGZhav7C5HvdqPlGa4duwysV92ZjEJihPPIBd7+3QL/F
B7m+Yaya8WUIrfFydB5esd1Q/hM3ct3WDet9fYe3tLifPpQT44SmkKmA9y714xJ4
D38gIDMzmYOsYWsnlHWilWmQRqg8InjD8SZhQwWbykzm2vISlekPLp5kZbPuylGN
fK1t4kvNTShpMyxKgu67hgNIm1lYdH/Hlo9sXjD69Srkv7U3DHUcamclzgIEyAGu
NdjQSrWuBNksKzbxcVWKGnT9baZMBz1rdkFiPvurWqLzLrorb5t2YL+bptVFSbh3
n3Pgfs2LAg2FBYZGFGr+/QcpQ3WaJncDO9+SoBbJph0EY9uAqXIvKPUlfWYZDs1A
SznfSu/vFl8NOl6nX7cbFNUgXtJXbfnd4MRTSIvHh8Hi7jaAUEvyIrTU5cPHLNP+
irt9F8wPt8p1XJo68GxWpgJh98/88gug/0FL4sMq09IgGD0pFcogYYPYVb72fqPq
eTNWWrSCDe1zRvCwTrgCy/8W8nLiIIw9ZlxdNYm/3muxvCCP4RvGZf9zD3oignAZ
6t3+NXOPBrrgzdcgc51TuQjgsO4qKZSYH9Kc5bCFA1DKA2AXSzuWZnbUJIJjQNvq
y7TITQq7npm2dicPpt4QoyB/6O49n7/w4cD+NwC5VzLWJsXcEQew9aK//ggYDzwW
Dfpq6XTPESCzhZm3ruN8bDdHTqn228lphXfWtBFIlA4Vy8+M4pkwI889P5T5+x+v
PolLE4ZO0GuHlvjSicmt/5xzDIWJF2WPex+BgD+F/0OoYnY1k5JfC1eqiHLAlANR
OFim37uCBfM89MDKf1Nc64WhnRf9mM01nYi4u885f2J0EsqFaGGPg7pTU+oc/X3f
PotjAi0epWl8CbdnY9NyU22ZI2UsJF+3gXMvmSVqv0VxB3VhZa12eaS9M1BA4kAL
Gtepmer3Dy37R5XZj+i0hMA1w2ufn+PQnsk+9pVZ4KwjR5NQzO8UZ9ZE7KpQR85s
Cb+SwDBzkGa46HSLnUaITZhKQfFnKFWvC/go70Q9tI5PwIwCDpgTb2Wi1KW9v733
v0JinRls85+P1wuMjrw6sF+HJoNNR5YUw1bHVPIMpRHYuTPAYAOML/WPNog23Iok
yDz4xLrFruAZO0Gn682523jHlhNO3O2n3xKM+KLGz8qQZkBPSlJwjWJpR+gqCMbf
lXgDaKp81ep9Lnr61jwqs5+44V5GBeM5K9csmxaZvMP0WEj/345FRWOTgsFpZkvJ
Cf6O7UNRIVPEziTpZz7HmwUrNuY9bnr2GSmweFC+BWH3b12EpVbrmozbEhvpUEb8
cLJnUPOO/HuVPHVgtanLEueKhODig77oWijComgdKH1NVgaakjtzcMfkG9US6KcD
RNAB+Ld4cgC8QzsaoYZUWm2YDRx1d/kl+ki9COMKRUOWWFQ6Zza8cknfOHD1rSFx
HoHXAGi6x0wAn9oNkVUtjX4jJI1mVHr15PfAHT3Wgu4i8yrzMOoOlG4d6sCjSCLj
+p1W38ip27xnhZv/Dk1jpruqSdnBR5M/ILypCJ0I8g/YHpO9vVvyCUgpH20cerw1
wD7zk/sqIPRkQ/GDaqlXQxWmCipEOOKnpAYmRUS+nt5RWN+zCVyT/4bgM+6sV1GQ
I7PMIDx6IR6jc2kHsEEpKE0dw+ZN6rONAetdVFFbC4ILh1gu5hrowO5eE3K0UkPn
9Qvg9kyFTfbQMp0fqVTA3xhFX801f04hiKoIXd0+ZlHZLEoFiiNeKSymLIf6bNH9
paRLyOYdDEhKdJpgdsPBAb+CMLLcRBs/BMHJkz34eihnmCb3LXsKfzAFjcnc+y5V
L1JQ3NA8CC0EAI9Bzfpp/jQNbu6+OFN/eUXE01nL3EzLhZuB2oWofDvYahni5HeS
jaV6oDt/tALp+a+3OJxcC0TcVsW7aHJwtszR+uRf3CLXBvvpSJM5fhUHaltmY7a0
Vsc3Q+7JV7+i7nhea6zPbv/3H11rFzDdsaw3iG3iq/jMHllVIzmphvdkQf3wlq0k
DuXW2Vu3IIoe7lHIUVafP4WJcLisqz1iGZA+Ktm2HkVcijavAAojPKVvHv7fHDUA
M2Sw3iwyS8dEfCHTOlcmDYnrJ0uKC9k/OxZEIvphKghwuorTrSSWgb5BM0LHPuCm
FhJpFLZL+cSbSWb3ivUTEt+U05/SRr+bkx4E+iCU3oZrT3OWzf36+FRfoZIPlr9P
P5ZYvIlNYFPDgM8O18AIMKeviHWTTVqwJK5pSr/5mDOtNdY/00JgpFCVmHpRhmAb
NVQO/95jhlb3fcdddQXF2SyZIRharX/Z4EtFMF0U15EeIIbBEMo8NEmg0u5Ggnm4
nHtelmHvCycrFU/E21oN7aFvrX75vO5SCNr16w+t/Wtk1QQMt2nFa5+VoEckEjMO
t95/0Y7oU+5hTdSfPGOGuvpO8uQCdP369PUWdPNhKHyYqZe3i20B/t1HCmPfc4mD
qo0xLcV3vbDuIhtSsavQScYVFSg0fYfgXANOd/zlSeiYcur+PwAvEntkjx82ZM2S
W+NJDyiGI0c+JCa54AlXAxzEotDqTU3nDSPUr1SGazhvoZDbevaFtuCTwqJV08ur
caMIRiglMR19kFNuCqadCg7+mzqawxDqXfLu2FIBUb+t/RsNOkw/JiQ1SUx1OB7O
ukSbJBkdc7qvUuoYPfsxL51jr8vsFrL/X7TVcY6nRLuhfTFAjQjdWfTyaTwzEU4f
ZR0MXfni6OKfl5smHipMC+ebW4cDi71VeCJeEGimAjGE+0bHQi0MxJL+v3Jflprh
eSyZ2s7NYC43Vaz4vM1ETRWCNlhINr8dDLolM+XFCoBwOFEBAD1L27m7wLutbomx
YRThNVadTzTABIk8aTOKkcxW8DKx47qsQKeRGLS610jU7nt5x01feLudSav5JBq4
dG2bTmBhih39W4nA0HRykM2FgB4O3LQHnhpRknpu6x9jkDXCOt8B8MC8/rMPCTlt
GGC4wy9jHpmbM+j0CqIvxhmLd/toMaXYFMDawZe7F/HsYQyQ/o5ZUqYCYBx4bTLM
BsVYTjrjCOYM54Xs75/G6g7dqHAvbWl9fknpH4OoFdQ+cffqC+wF2VGt+mUucaTQ
jG38zLp9oCko5FIVaLqSpKIfuGZI3WJNFl+YFNn9tz2s3J2639vFIMeP9tc/jisD
2ZVTtDW3+Pqz2cjIagqFdnGLNB0RYfYcnOL68ihOPtlVIo5a4WuEZqXdSZcCDgUV
gl/2t7VABwMEr2fVOcc92CYgu1qV5sS0mAULO+TKxR3iboO/BXrWKW60oOsKmB/z
8B4/PdCAudE7hcJiqZPbKUOekWAjEBuZtFDm60soiCiYUp0WpWd487lt5sL2Bxcv
n1weajdlPf5C3LZYxKlXcKOoo2dqWy1ZexPoMcvqDBUljni1esEIZuxpxWwVIHsS
n9jpqxRFmxYdiJSAeoq6mNmzzGLAQC9PAp2WtFWP5okFd4zYxBqnZDPJL4kjaKTx
Z++3CL7/H5PNDdIHmSELhMi4qYSWIepv4XBv2k9oNVxGTKgt/+UNCJybX9a2XPBi
Cca3pZKGh05surJy4EJcnyY/ZW6Afcw5WOvEyj15i3LXEExh5B+8OFKthTzk7U42
M5MhzEnkva5yR3TnZBJLABQv27wEQQFR0JASrzCOW5VtrsTE3yLO8ib9oshYis3u
I1OD+NZvw9lg2X1LEK7JimTIeF0ZitByY5F5O2JNsIUKCknm25f7YCC+lTxb0Nhw
9iFAISS3q00WN+7IqHyr9DIanrkiJRhITQr00aKv+h+LzNU0Xu9uW8IPOdcZt3u5
HV0+JPe3GnuMhscHtMCkZrGKJp031VueFW69YztzhrmXTHocDf3eFt6fOcregXsc
zPvAIBFaoc1dPXWsgEmQYdz78ER0RAoVy5MyBjI2ETDQTR7rXcW1UZ/yrvJhdhVd
xjSw0reC8Ra9Yb/XHgjNBKiKUggss+PuDeVcIe88M49Rve3xoeL+QwqULSR7EBs9
yV5z6yTGLCWGyyEDJTBnVPxXgLxU6O1YmRBxGLDJIEswZ5iVp49oINA8TiVOh/c6
BXW5UWpLnBKgjfzeCmV4kZtLKgi1u51uNcgKMfd0GT2bN1a6YGW2m/eDGAO/OiOp
BJ42UNKF89mEMH0L8Js/aVCN0aA8OH3LGoaRMpN+WCJydV+LMLPDan8PqJC3wf1f
o5+ldY8C5DyXEbV/WN5TXGPyslpdeFN6Hw3hVPvG6+nEG4g2tg2Zltn4EjUExwE1
pSpzLm/EFYdDZPZIjYfwOMvM8ovX3Vr6zGV1+M6JHUuiKR0NyGXDAS+FhFCRmrxv
Wb5AZ5714hSp2siVFU5Bs/VrsiyqLTqsPwQ5QqL2FYzMHC85DT4YlhQ3ev7VJI1L
sQpxL0HDbKN/DDEGUM5xbTo4xKaP79ObGtlORLfY6Jb4EoxTX85U/CA/SiPQW5ON
yYwxfTWxBkfpCbdfujIZiDk2aQ9njfI9gDD7rRCbq6mg1kj21xLz9B2MQbnm8Ms9
8+x8ORBBd5tkGn7hfyXFLIEl6pyyVAzu5+ea9KnnarpwoGK8C39EQyMUR52z0oCz
GpCVoTO69CLWLP+Qezvbm8m6kT/NVoeMdRJooll61DILpBnRi+lpWOvL+OCvZvta
Uabox7FG0Z6syM0MwcInAS6cSPblNfzh5nPpUKTQzU7fsySCpbcCPIb0JgS6qAV4
IjqTGt5otdjDlgXEzmfx1W0cR3z04Ag6e13UNLsWMeU/PN64ioptLPx5JveLOKdC
GUnCPkMb730zpW87UzvgoWvdR/FULMbBJP/ckBcpIC+DHd9vHSlU3YvEpsWqze9P
2Gd4XqihlVBZf5VC3ZiY71UfrQ5Rx9zIcYoma6j/p54iIiq1zlOonggpjMDwJYS8
RbQJhHo1BDHCgVD8g1/txnJfpGVumO16ibj+x5oU5UBtU370s4gpUsNpOS04TR9y
ST1C0ymYZnm/7EBMVbB135BysbvBHCo3YrcnI+B/jnRjxnaVKPsryyq6ZnWNafcA
hu/+XpUp+GbP7BMOAYCn+TgNN/n0B2YYVQ4ODw8kpu3AmtPYucUbJCPAkPnwQMu7
hnDVln87cZR7omueSThHT4WuEJd7H7VqyPfOdRYDR3wcaMIBemyDBSnHtHMJSYCD
7SsK9ko5Z2KVShaIcpWTi8cIvAZGkGVxBPS8d72H7EiCtRBWge6CIOyZKqu10ZPK
sB92v1cTCZCauox86gczi+IZU7kPSlayCE0xCqxmsY/rjOzDktHGSiectokMv5xA
mnsM3X95PJTo2BcRJY8fwExiTtaHfPUiWdKoa01bUn25eMBcI8H7EhycH0xxpQGS
85Od1OeXeLCNimNtQjtJYg9IG1JeyrNtSdIZQam0woXJX5O+/GVoJ3IZdn8MvhTr
zVRsLhnW90QHc/Kgme8+U4VFmfNSdyCyzOGruCrjL7sqlfbuxkH/XdznDpFCTLJD
qYHF19lVT21lzmB35sEnNzbzfZzqHaWuGZQsmI4Zi5GcpLOk0X2ky8vSva/CaS2I
ZArQn8JupRUgVGO55+Grusbj/r8T3qDCYz5xDIkubKuVR3CCAfIaxk23tbevipiE
zUZIGetpiLIyI0MvmLYCQR6oPrcFcQtFfNO6818c/kGhtxu3ZuLLENIWOIzMFTAu
oOPfLcYaZr9HZfjtCs/VakZMujq9++gR3gRaObm8rstGc/YKooME29HF0uY5PVw5
mmbNF/whGyF6GtZrr7gcASYJLSjlkhabJWy61tk+U1WPQyycdlfCKcIsEprKqIJw
9gEG254KjKCqm4SjHwBjVXaLDks4FNuKKByVf/FFm9pTp8SI1yWPt3ljWfDcJc9L
Rhy3JjZZxowOEBNXefeYS3jlj/AsYcuDgCeNdyIFYaWacriyh07rb4affSpVtxYB
ozKtZXnEzMFc90oLspv9wyl73TXUtmCXRvJCTAEWfnD6b1B0Jr//KtNkL3682F90
7rGchy8DI2KycIUe+pi7e0KHNhjPUu26YI0XPjm5OIInCWKIsCOfQaBE7XxeMlYS
UywruovULByy63HJpavjP4urJvYynwLiwmeDICl6xijxtGFCmSGbAFHCYC9D6jeH
cVc3H8967K9Mtcd16hWm0tyFSBNvugA2er6iuQSuk3+3DUMfp5wd8S/2N8Eq8uj8
ZyCgSURhyto6pm5lKMwcP3x5HJ99onCAsntbQ1gAtDL0M8l9UB6mhVd0rclW4KEa
YlaG1p5C8q4Llzulfe9CopJaPs7Dc60KYxiNfTVmuZBttRUKyRhXKLn1BQ21aW5Y
WrYQTVp+JlyeZuEtaOLI1bd7wd1GOk6JRrOpTqoMJmnilyTTACPl088io5w+eDvj
dsnlDQTNVn2KtW7wU4YOYq1FxP8LjelB41zGAjjh//xMB/XwPok5Qk/QbkDkkC/8
iBN+3aWsvYgZmrSb2LvWF7Z5l+c8uQ3wv7RDhTSGnhaGds62PQdt2yFUPMv87RyV
fvujAwWkTh/7I1zGpPm/p7aGxgVJJ6/rjrafbX5Oh6lbMWvbYCZ7tIvAiwMQsosg
0maVeL9rRAGXOgwvurcOcl3uWRrTkeLUQs+JcvepRXcEfeOd40LyQDIlBNpSF7DZ
aZicHeuEiHHHJL2wkl5qfVyOSmkcPviGXiOyAc7UnOTDnfGAfm/XNcJPE/GNsEfJ
157nVurdHbr+do2AWgyURJnULgbJOWg+GBSfFZs7ycw5oMFmNNwANPLyWpxfqAUE
m/XV+Y8OIowyHv4NswtmshI5nnUwhpcKSYrtPCpy98ZwFmSVRRQf2toaAXnTxFXj
ppWukuxB5phPZR67fywrJllLsx/ckR1r3e9eKvqi3lpXAM7dia93byGXIN+MSuLc
315d+su/Q9D84OZoeeUjwpHpoZl2HyAvTeRHR4aDEyzoTVc8sNo2Ell2Dm2V8ovh
lDbhVvy8Suk0Lz1dFB5JPE1OIQMJpu7qnJA4uWSIi+RrFk7BDzQJ7o+cC5SCgg7j
XBhne/YVK+KqYQftnSwT5nRlIaUF9tzdS/s1im7YvGG5jxwAjwAjXMA1TI5/7h5P
+nO+9NUl0lRnR9GfCzntBgXeXpo5tWDth6ZwtexePeTynuHWke7xrc5If6s1LEIh
K7Zqz5Iqt97k1k1U1qE9QeBMsUgRk5TopVgFq7SACQgYNaS7qVlYO8UmRdzxEJcl
upAUdxZc/+N2IDGTpkGXnvdx1dDqk/7lLeUZEgrHJx9Hnkh+7ZEKIyGCQh8Wcqno
2SD4C7L0Jf5bQvbxXGkMgBiITYrrWC8yVzwyJIk5ikNRQkPIqxrZt8I5YuGrp5/P
2DDFmxUkEGSEerWCEvcyrYLlYZa2l3tCSnMTVdE+BCIsAP8RFdYAZfT+BAJKkYk8
T2/sOxkh0xcQ4g7pHFByodIHwrMPBii8z9BG8gA1b6x3jyUv5dQGmG9cgoTLXXvx
7XV9XCNuBNN2eHhcMFlklxrcgtx8Ht3VW4TsMYedCCYjpnr51JWVUSpYFm56NBlP
5dOAqHk+yxNXh2mdox+A6OSo6fKEpiu1jhi95aDwfjh+Fla9xKY0zADgksHWIpZu
pLKq07LmIlIQBgJaO/cwVi4I0XGQoNDQwEQcrElZLVIGDEHyU0ryShk3erorBqh1
NusloL0tn/tDej6dwNfXrYrmFpn2IuyZksy9G1gfrV03CB/2DcqqzbkoO/3dcloR
WVKXVaj1qjrJUKM9JCupeCTvepswTzQ6mEIkcD/zsbMX4SpoqpTGVUQ2AxKlPjto
+K3P6KXnPrCwVjlzNT7GTQ6lmE46UUmdMRS7GlGRIBLYE6kNYehfOaWlGykvstlF
kNP3VSIM0tcwitniNFeNGMmbHDe+upjb4jWvHazuhs57BwrgC8r50rH911YypT5a
6Q1tfz1EvzLVGpk18IX7uqi/7Wck+KQL1ew++Lk5tcaOF2VVFZU1fqHzlALWTafq
gmIlqLYAXCf95ljUvcIR2Qzbful5nL9heIUBSesMXxcPvzlg/KROp+tJemuWEg/F
0GOvq6OrlSu622FP4SjG5cTsOrcIBwoeDwuwq2dd3MCziEHF0p4wsUMU8uipfts2
Pz+CnpLATxI3p+qY7owQTQ6485DBfqNtJ23ePibJp0K/LQWiIXLgq8YxaZE2NYp6
wrqyQ5E3aJCV/IHlf4cvxnpHB9MW/wWcNzk7SdQw1O4p7v2mBpccXMAKzyqgZenm
/6a25csaPCq5heFzHaU+3Ip3592FIVl1n6VG6wNYmbCq+kJxHNqjnoH6yRToRlYz
biG1tkXayoWoKjeDyJmjif83W+UkgO8i3v6+NASFGNmBWY2iTHPme8z+GgSXKnkF
z2ASZgWWBmrEXGu/Y/UmGW37mzU5h1FhY9XiTwJsdF+RuTHa9v0OGt5u3ehRc7/j
rBS66snH00gNPxWWo/JIRksT6QrUWI+oGi2ISylPqOEbFCyiKgxG+tPo33OszCph
ToP7DMZpv3YZxBVKpMiqIK8xQlgCak3yuynp+5o1EngRWyma2NbY0qkHMeavuXFS
0F6JwYCVuEDZT3cM6NIQnxRZiBJdewYbgDJkDpnRRKR18snLpLD8t6x/U8nNUJdC
WgjalIcZ/Epo803yi/u4lmo34kSbIOMowz/J78QHYquefth2RhPniCeEKkjEO/md
0j5JUIkgAvbNjOlI3KAjyx551C9CsvxmVr452nFg5pCVFcVoCE3slcv1XMGfCqBx
ohQ5i8P5sthA0JtZz7MblXkfmFaemgBLe+kHVqTx8KM3ZVBuh3fLsde8J3wt0Dk4
/kTrsmmble2LJsZQ9thJrI2kt7HpgnwDNoypFqaI+mgTEu+HwfUi1jbRxukuvUK5
jfXEN3uYGIDcEwbyDIlFTIel3e6k/xschTX7Y5OUL3Tt9JocrFduLx5O7j2R5r28
cLkHwrGCemZj7z/cDDu4MmB1ypU2auvwQmUjLu1Yg9iJ92l8+oopbn+D7Efz4Ufm
C5JB6yOvevfwSW8Vs0SnXs2W9ENvXGc+rwBOyIpcykU/kOVvxlfUk7MJBnagJvQt
FB8LGRsWZF/AfVJlKK6xLQDptkCUzDssGxORe4cBzwEa4PW+c8JmZsqyongkoHDA
K2cmcZAEcbCVIZ8YTcXvThnND9JhJklWv9zlyrFjTsXD2wyjj0ftPAHWNhGjYWcq
hwwB13AqVDERSs/ZYQTuOryIxfUd4xygzVuBQz2BRTnzzhAa6fIHJTprXc9KR1fi
wOv2fXF4PMyL+lsw5zW492it7u6UjSboyQenloRFL2eWKElOszz+vVsB0HpgGqNg
TuZMhPdHyHhSsMAimloQAG3GuBnwOAwE72MuiuKp078bLUgi977p5WTDEZv2k4pg
LiJJZ2T1reRsFVFsvtEtEx7SJsuj0qQOdrXi9i3ZNTOwzdrMdJaOXsJ9IzzJ9h1N
FBJL5oEmrKVPOoABlQ71E+p/MRIEU98smTGV1XySHc8HtQdlbeejuTVxrq+/1qpA
Uq36dgZlvgk2qh5TPKEtKCzuFRtZ77vw7Q4ORwKOZILPxkuLjuyYGPOufig+kgXk
DR4Hrt8VfbsnzemRKl05EdW4pkw1fScDCoJDkYuh4Uls92ePLdMts85oYy8vN6VT
RatYyqBa7FveE+zWR19Z9FR/3QVr9veJXbqnUkusnA8Q2A/JUSo6NFssFr9wCbQN
BIYlU2Z9fzDSPgQhb1f/Ti39G7j0qp6NLvvQb7o3EfwwfytLlhfDTkhIUfTmxrr0
40M33E6BAqz9PlWcC+xlv7eiA1nxXNLb0CSkFl8Mk/wBkTIIey3WMHoHtbeI7V0I
zXZmYiO/vMiVFGhy/4Qi8NxSj498d1K8N9Dv/6ny5l490qgxvUCC3P5Ro36ty+HY
cfeo4NvIuYcfS9fhB2RTFAztCYFZUjxV/nS8Gnr/Lh8WiAheWvbkNfC3WaKwc4J4
oFlXDxWEwGKasq1cYkkkG8zCIr2zg1t4l0WxeMdeBhyEfSzYLYNr/bwuUKS3IqIu
J3ftELCrc+PSLB4oXOeVL+sUgtZlNFoocsANwyKGpwV1ji2OmOxutMIpUrfdKCj8
GVGuHGV0xO+fBR2iYOLg42UGdBAA4kv4/01S7fKLn2c4VY1AQo/VaX+dcveZmpOG
5N4HYZNVHe3Fnvo1oWHP9dp7NspRqS+45y3XSnPNhYHtHMOv/bmtR9fbMeU+huc5
3LAjNgflvVy0FuFbD54zMzm7zDdLTySA6l73d8tkoMk=
`pragma protect end_protected
