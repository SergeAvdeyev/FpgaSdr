-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
b8tArWpmDzEdydNvlmCT8U43XcOl/e/PdqIcXyWcXhcEM8lRc50pqxhPWrOf8WxQiB8ZKvRaO167
EgGIn79igYB/IXc0eR63unLK59UaxXefr8+37EUBQyo11LrjfROmpNUmYSMucKrwqem2M0cop8JW
YlaGpuDJYfGrbWpoJhpineRdM5fw2ieAwBBEf6Cc0vT7bzW7HF63l3zYPAkC6OTt1274pFprgXoH
zCC/BDqiFB/1bP8jakOFu7jJA/yD1SlzEz+dMj5ODnj0YI+q0cxsa/B+RyJv1YiT0kA+hyCf9/Vo
r6q+9xWNb3S7i11+Ez7sHpVTt5KMkUfeXWfRFg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
EgHuYNX7iIT68PwbJ5C+RBEsBUotvstmZSwHyBLG1MmCSvmkWdXyrxGIm6d12UnquQd+SDxHL2hp
86vHyNE4wqRFiU/8eG/eyuiLulg+6cpY4VhoA2ePCfoKxt7kwFZnERPYXwZChJARS4KsfS1XlIfj
EH6fQihF3FBYueY7VBRCMCbv+RMTWIHiE8B/Ihqx1I5BBwtFi9umK5E9/DBdtpUt+LMTck6MuC+D
IFypxBKokBfWNvTg2XawWAqn3SCrW+9c8wnF2siU8GPd80EuABTVMoY6Ry2/kg0DV195xIO+rHAa
K/F/dQSW0FzVqdQTRyjY1dvJRZzqh8Nof4OHpGjc+rRi4jATbklnq4d9ds11aNGiMlRBTGIf/seO
a9tmwEmv8oVVqXgQiVvJFWETLybORwLlRymla7QjPXRmqrRJhA66Pbp9ouPte8TBIQoF78z+myUJ
lU7CIBo+3ENhIaVukAAc22UvlK4rJGvXlCJ2Q1vKOPF+Y1i7Y4r927D8KwUSWCB0jagpToVqvEIn
1CnYlikYAIo+8r9TFwvac+ZQgmsLsqDu0JnCnbjqMD5mS096FlKuw9u8hkzX10WMbniLPeqNy2Yl
6EyZqTIBPV6UkFsETp9scoEkWc2S09IT8ZUEJzsN9d+1scPicq3f+SZlT+umUFMlSOo4Ktak4sfl
40Sqy15iqx94RTZaa416FnLd8Pz1O4ohTeOB140pksFVmhlIXYlG4IDQHG5/rrVJzPY955sbTb8v
Wk/MBBBGWwjnjU0lhRaSCVd9DiYrZY87WCSzInws67KC/lNQ+NDpX+5NoK7vvFNP+IdgcZ3EWqDN
CohL0WgtFfqHFq85YanKftzInggjbfkuftFMYD6H3LFdgtV7wIBqU4hpX3jAWbBv4T/+27QM1iFX
9SUoCS8Qtm5+eChIsNXB5+q3ESHVyOt5WlFgTN3gIX4jqpuGbIKZ/77WOrfeBBVErCtdtwLAgtFe
SO4q6v7vPCYsQ21PcY6SWAPZ+qCR4U6PH3ru6+WdYhUlAm0vPUxLM1iMiDT2gIYLR9lnEqemfHk4
zZM+ytEFnl9mwhcgfmfDDyj2HsNHBhGThlzWYM+vPIwGB4bn5Uj5xKAhBkPJi1x2dvz45U3JXvAZ
EAWr1xvK2JX2+57Ja32vWR6hrzod4Kie5uaeyNuJoSX4u6pEFhqDZo+xtULZtcjhSEi0px18YSbt
8d97Jt9eXh4qxpC3CKrbtOihGNtNpUlcfgT2icNmKVWX19zUzxEqWv5PVQrgOVsbpt1ds/FozUf+
lyGGffQAxF07/GVRgMBhc5zhCS/NuXs+1wy06SI0NTP4bY3TKVOhMEyrdVr3JPf6zLivdWW+5bRD
z/miiHXxzEH9kYFK5Jfw2/Vb9B4vLwDdxp6OIL+4aBkn3IKjBImzRfRPtfO7U/YTLjs5RVrYBKmR
Z0GuuZHR7TiWI4wF9oLy8dZC2Gf08OvDXoQ4Y5AO29lIMP5LOy+vpjSsMlqSoXR4MmseEgPQuL6d
YpIzEDhXudoiDcKqe9G8QYYipSqMIdG0OX2c885Q8vAtbUEKig4VfEBN6KqX9AAZwP7sdTEPn8Ca
NSj8LGp4Kw/LrUXFtubDjDFdK+5APXaof/kYLLG6GGLx32eN67v1ZmTU4BNPvsBkw8AWulSO5QK5
LVAgL49o2rwsXnECoHowTcpAIdDEdshVKeNc/Gj8i862G9QXL+aUSD4W9yvQEthM459H2r1x+XMM
fKaou4OBSuwAknMRxIsqJTXcw1VtwVn1JgG7d1LIGvSsWEEQ4zxjBJe9SI1Jws24dxQa6QZjyZi2
W7F3CBr0ZBFHQ+DBDkGYBXVA/QS4LXWRFpviOUYxC6VX6KzQZB84HtIucPXS248O0aAz7r+IR4+y
2lLVSnvFanpKjdJbX4IusrHrpaITPfnSX7Y9fnbWW5vCHKho+TsMipOUZnMep7R+L73NBkmtwRPa
llQ77IKWoX1CiW1TKpoXsBAIE+he/6f8l1GktoG7UBwMski4vBVBJnOgX/h7aOlGUh0Hhs0lFe+j
pBry7X+kkRMOucdPTUkLHTnyF41Vk5YxBw08nFiCKnWRt4IAegxOYoOx4E53Wy7HriXyGpuVSj0S
KiOcb0R622y0BKUzMYQeWxWDIIgz8Tt0F+AkAlqS+fHp9YqjIKY+FpjV/gIPIpsFLTDwoq8mGJcr
9FhQG6D1h0pT9RHoqsjj9W9HpZMrPknzk1nDG/h9WpjovBZrIg8g3Rr3yx8SJPYy/mNxCsQZCdUn
H4rXz6y0UHCgjCHmKZReC9BOp1vi9XnSOmVBIMLSewEh6whSGY1JPPdQ93SklJVkjAHsfPpcBIZi
P3hqz53vVJkx8KpnY/OVfs3p0+Ayu0U1QqlCJkITVOsvlXlOhltpd6ve29CAWiPSeuaJII155ngW
thUjuL+1xz2A/nIrwRfKVOA4ApFxoJ5FGgyPbofTF3r+HVibqLQoxTZGSYINiS9kh5xnkbT1u/Yy
/7NhfiOsCsDR+4I2c4Q9ZT2UsFlLMEdy3+f6/AAYpDj+/fFqUpAdBQEpodR/v8iQmXDBiaMAFU9V
XyGrkOWDuke4sxFMCEuloROnPdhBqzjbsoKGfC7a0Sm916OJNMdF1X9JEMtI7vJQn3KtWiSTd0fK
oss4ObGtrBXF6YCLZk3Js4/ZYBSZknccHSwHI/Y1fqwjwX8N3DTgsPt2LajvMiRwKCbDxCRRl674
2ZCjPmWps1fW49KLool7MKmIf9nWT15UEYp+nIKnKtqH9K26K4755LAFEQoK0BdhwhPlU6ARk3JC
3xcJolLL7vllfXdAVRu7IRTSnCAGcETrObrqa+jhdZlJ42OeTk8pnZ4GFfxY2Lwa8pSkQF4r7CEb
LELcK4CJyjisaPeXgZSAgsw8PDZNyeEr4WkDTDdqlTtYlN0dTftQFlXsAQeyU/N0GgSinfBWOSUM
z/5BHSya6jNDnxGBYbJ7eYiM8lNbCKmQxsMBubQrV8JmR2qvldMlauDRqM/f5pXNpkACZ9RftY5z
fTxzVKdi7f0IrP52cdpLb2wVrs/rUHyhL3ufYMn5UohAMY5qxNnmFM85wBVyLtHh9GF/+UHft4OH
jQ+DE5+SgxXs/CJQrXXyO2o48BrHdNdAWw1a9JoJ+Q6d79415QJ2YA1LZy9i43hQYYaROX1P7a60
LORfVgNuM5ICZf2kDDxWdeVEzrKgQiOeZJi5Q+VzSBAvuueevdUVAK3XT4fdBAzo+/Ke6WSDYIZU
UIyMTsylnjGqwtOJ88DD2LHJWDDUJ6JQBUqXJiSKB3Nio8wOQyLujrIfRup4iEWREF9DZLa5a/fN
NAU/MZtrWeoLcbeJGEV/FMh6jfacDWh0IvjF/Y05u8STMh/ciSZfZyqFeLTTBTLG330HWnHRGtW+
ZUFHzrPO4WURiT8dkuXc5bFiUEcTdPncdMqUxXTktrhODGN37fb4+CFAryIcE9P3pRoX94Ab2CgP
Yfc6b99u2JVA9VFOmA2r2NrOif3ZGHN7/e6wwUy5oqzfe60Mejyv9X97dOT+E4DBZAwS28IAqHNI
TdpMUUNrR/D7LXkjRwQG52tiH7xJj/ee+NYXipQcPp8ahAlVnVB+ssLu7ECSHYMRPOf60ELuKeUR
UwjzExB3GOoAnV4QNWioRzAwlrcAH6eIWH571ehq0hTHmdgE1mLopzEgM/m3k3jkSSgLdCCIigdy
PY8N2dEe1gWZW5OTI1Hq1LVxfTY++1mp9C0na8KmiGj8C7TCmDMHsdjYJFFVYAQXfhvFd4DoSzN/
es3/sXGDuY1HzVL5s7sHNBn3C7ipiGJoJHIhmCOMgFHxfJvs3HgymmZQszj1cI3TIjlC696cUISa
+ayFHn+hPQmUvj1Ii5pPI/W8yahhu0YFGteWUIuddm63/dx+axQ8L20uCvmak0PavM8Q5CscxQSY
zAue0bN3HNhPGVmmnDnqYOTWBIJQ2D35cZXLssPsYeV8pQJoj3WY3GAbiYr+yWesmOgXhrwo7dC2
1pf5s8vX4A5iwyVmCPDd113ijIigrQ7m0XDu91HrhPZrA32uPdcTxtDoEIPMoc4lLDJuqAcFBh9A
e5EY+nH9xiqI0tSpO8hdJOv1PfTn1wYZnHC/mzMEKp3qig3Hce5w85QcJlPerMRDIhXqeCwxzeiy
pUIZyZofodHr43QHVhjY8YIJdvhdDmJg05KzlbJk/QSS1AAkNTpNWJF2LU9uDv0ImVboZ3kuZejI
Q3ayjBTvKLUGsSEMQR9Gpto8b2hajUInQbY3+C9+JgcaIunoHDJHCWEOh/ypsM73Cp9/84+RVRbQ
uPTqjDcBz9mPTkYK4mXgPmNIz+4mJu8+LmbQIToPcDmT3t9XFMvIaId7a1aqVipDv6zabm7FubxP
KIEtYV/DRxDtzGwv0LkytkffB3F4wMPj8SRGoITrZBXJyO6gaDGphc5wAG/ygeklmvg19niUwv3D
GZBXDQ1hJdDXE4RVwQ0nwQdloXuYXzHBrpP7YwChMY/vgb3IdiVmxRcXLe66kgaTE1HN+cZ7MKE0
0WzPW8OYZJ2HFqz4DqPtDh0vAAic3T5TH18vf/4jLQvDV9UsbTd+7GZgRpSm/NJtzvaDeccah/3t
LDCOk2j0BSL3W9TTKBbyuFia7/Kr/Sjml+E5peumtR87G2O42vs622/o7I+D1J9b6MkJg/QP4IHY
jSV8wUi42ySQMZRK9LOPr3QY8bAd2ND6TCQmKAeYkZFyjddKTI6WQS/hGnpKLCDqeqeuWDIGC3wi
5L6QEjnEnQklel2a2DICwyYsMJlbzbsWdEr97fW9u9pA3Loqf18IWvOvOwuSwK70VdnYrR6vZb32
14r5BlTm/5lTPMx/YPvmVStTAq5vMcbhCGfJ9MLwXv5N5pGULa0DFcEy7N3NyZGXFJzO7HiqKDh5
GVcLEpPeOvZG0LBtd6dyCKjskcGCqa1s19A/ENAvnAXNPYMpP6sv74s92NvrMtXpCxaJk5899N9X
pkrWJ0bqcqFDJsIkyQGbfD7ojOhBDl6V8gcv0+4Teb7bwxXIPW71cKxHhTdG66dzUbOFRMnbOhqP
xq+zmPmFsMkjkCLZCy1vyuKz1OSDR4yWHHKqJmtGd9mycOSxgqkCzlBPa/BTv8fUp8B6VeWUoHRx
9UJmNGUfqI6pXhQNmIccs7STIAwUOMi3FfKUQnDYRegJ4JX1WXYD3pG3qgeXpgmZ/fh+r2SgT7Fv
yFnO7fIMYE4LC8/OF/cDspOoFRPaepdI9UY98ijUFsZZocoltZXh1sSIlAEJq6/pD/cQ+nIV/+Cq
mejHfMz0pt2CUS38GKOHbWxYiKLZJnxz3waifDnM6BC/KzrCU9I3xL3/IvI5A4GMPvJSVh8yhEEu
d7CAmzdFU6icZnqLuYiBnXPzqEjJuikX0JzKf0SJnZnW98PsPUqlSPST2fD1u4cmoajcCO4z8NGI
u7XcBd6Fj8MiUfEvT2VzGnOdDKmjA2B5s9+rmdetOB0rz/FWIeu/u8E48qEZdQBmw6T73n19z8gF
icNekimZDW29fZAoAyJpTpx+S8LX6ZfsbkCihcY0qfo0XR9MTspf3AzEMXq/nluqUNFM8wPmsF8H
6rWlA0SaH+js5MCw6MKaXh25Ki6iukwDEV7R0Z7rAE6lXkNKdhUMjH8bIbnbiQ5CEdOQ/Fw0Ikkx
pb4m23OEb6l5BUwZ5cJtltePH4+py5mlhhr8+/DRNki/2IiBceRpJVCf1kD89k7AzjQQJm0MMooz
5ySXb98ftROLcuyMaAjb7Hci75TPsjrEFQL8GIf49hsmcdqhlb4SyzOFSg4szTkz6/3X7Jqun57j
eIecqJXYXgytEcqBbYW0T/LZTlQ+XHZ6kv3om/tI5VJKJiGnM5Xe45sUVrgjV+o+i/1E8ZprIl0S
xF9LhhBth0Sgeq8E29exAlTQSHwYuxEveVOVSwCeP1ZNWkFakS46ayJqQf6BgSP/w26XFpe/tHAm
OnYbm+jPGDWm+SiuYUcSEOUP/v4692cDi4obrw+p6vOyFyQPQZlWKkIYlGFc8yGKrPuj7r8xfhbC
+kYbxOoKScISxuyo/nm+pQko2ZAxS5zRFpcYwv4N0inWzXkIrJUuMjBxUt5q5MnIpDCVgH/SYEEc
deA/FZoVKCTGMc4aoJKBNDxkS95ZcXC5lXkG8wKk4KTe/HqH47HdM85OlIlnn1uYXPuh8dALHjZO
6DDK12v9+VhgnUILtWexdvY68T2lMj2B7ZGlaaYSlFNjkc456rNlOVU4RTBlCfIuxFiyE5wKuQg4
u3ZMpP013t1dB/B7GFn8O4fm+hx46XmFQpGAmXQNU38SY4s0+Jocy9pfr9FYEVWTMvkXJsf+W7nv
NhTKtFzpqaTMVi46DyYgPURrVjaG6+yutXGupPhAREeEdMGK97UQgaeqea3J6/4t/gswcD5iW/sX
OHzoItP9mjmb3QX846eG/ju0mT5rDy5bUOZZAesGFk7N3Mi2T6UxFB/fJJEDCw+JL2WhMAsfxOdy
yDi3ixQ1v8SzjkuJUk/x0LLzhmF31+k910s915DiAW2cNI1xI0GQczzQvtZDW9k2sPrhtUodrPmd
eQZT8j9T2KDw7YH47KTQacgMj9D+0SUKBjyGCgOxd03GNCLe9sG5XER5xTnSUqrsA+a6XLMYlBiH
TEiarKC/c5o0rIuDjT4+JnSRvowx/aA420u2JaCntzrC72fqkIpkF0fbqcnNzJ7coswX4D8e107z
DDuWrb5ewl1BkLLdmnuM7qSLLgtjhbmrxiyiIfBkdwtPi7q/xU12xBBFiI7cidayof5iYxgnXtPA
gpUcTOJS4NbbmGxsVu5mrS6lHAS6Nx4+TJ72p52Rpv6MW4F2GxWVAZuckRUSZ9hK+8THC+u99mxh
LBlxEAiaO3zybrs2kc3RgQuUa+TjR1A0AjjEwKNY0lmg2+TGuk0gR3E4gAmxgouoG5BJL38ZgsRI
FPG/umhO5V+SxEcanEBkxsedE82BHL571vFk5xJEe1j3iWwGGMxa+1F9mMbAcrIfZ7Vx41H0xzhj
0iWTOueCLY4rFt/lsoYVI0lfSjFMHzfdvo5p
`protect end_protected
