// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.1std
// ALTERA_TIMESTAMP:Fri Oct 27 04:12:52 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d4fmTyIrgQiyM4ymWMtTeYwhgRzGUeaQoX4wl/voYzIOOB8nyj67gAZMkHmSeCkH
07mIyP+4e0gJSH2tqVg6Ek6cQDk8aYeFVNZaFAtPQwZ9pjZAXtnvYtsQWYMmzZqx
nvYaDZv2tH/cqygf3W0i66PSoWdynQ9NSDa3QHQTtB4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
Sr//jCIoeEhbv1hLK0uyzuyXH8t//U0KLtjAsJUz9eP6zUme5IBezlarljs/Dryb
BXUoytTQ2enVQcPSG/otSg48Rm50lhc8Hu4GVTtpyXb/Vii51EHAup4VZfzg7d9N
SfswmDK7fJN6FV+F5NcyY7KlvdgGuIsrgCCSvrixo+aeqFRV69z+nbvtC+ghjQiC
SqGJj0ZFA+jASKgq7bZkW7w+os/zKj2yDnX7pG4jBbKfW/Er3XTSBcGJATdhxnej
NTsV1rnVde7lAvj8vAVMW7x3/9IzQy5ujnV6o1PtG5BYu+sw/3zIszANBEHUWEMK
xXwAbIhjiEkQSq2JKZG3wVIrwnk3HhCBnQXh2SY2y9Q8b/pjb7ecZhSviO0ALeE5
hNWyuxpW9JQEi/ykCNIRBkDOaGpYF57AOSQ+dbSmcz7s3FcRcLBaY6mk2ESqzb76
Oya0zvdqseUIsCkSFpnjArNN0xz9C4upmgJkUdLT6oZZ0wGFlkfUj+ax0odfsyrL
4cI3opijbUvinso1mPQHXE8PQV8GbsGHdQxhj3K9BWuTVp7XxSwKY435jTFk/x5R
vT9jNfqMjWA3YW7N1RrGadEzx9ZQjHg2FuCeoIeem8+tW+q5dpfIboV81fPzvz5S
JEYFrD2h3/X2MMTPecg61KxcJNrwTEYx0xWwzYIS6Bc6T6nrU1vQHsHQFUFtyfk/
6VxRMpXHxs2jAyjFbW7LYRiFWagnmX8Mo+Nhkba9mShNtpJXShEF6deW+fEd3Z3A
3xdMUIta7BEX3zMGHAOdROKwS8oYQL0rYFaQcfB0MX+8Yqg1Z7h8v++wLmDJ8dtc
3+pm9cZpTXIoLhpnvi/wvObRD02xpRb6FkvGMitPsfYkxEPKwWFn057sVtDR5AIO
BzM6zFjAhREw0IIZOM9wGDoV1OyFSRe4naP/UBDIoAcOj+Ii25yKVSEalyAJmxBc
xWtHin3gHnvXftuJDkE47F5ZfDkdIbZHFMh8s+L1+RaoA8zyPiI61Q5eCH6ZZkdJ
eV7P/+7YM0Gv7a0EJIpqeCia+wdhvPEhZ/1cKDsQydpe58rPUt7pIsBdQmAf1K4H
AxFrVuBfxEOm/upv7m51XlT9b3yhiJoWuFwjl/flu2yqEeDy6QglUlcltcuMneAT
NRDnzFTd/CnBSriZljgkDPPK1vPQ3uMosUkBllKSor64RPheeMMXzu7iRJxghDth
qiwo83TD/kq8FC99gZ2Sp330eqt3OlDXBr5vS3+ZqIMoIhmjq5JH+bHnAJTzDkPW
PgA4G2fBZTJresP1LVSyaDWk6YZamw5drQEmYbhljs/A/t/CEp2wIhUI0v4QKvc3
xdSEV0yeT+buf0VShbYzL+JfUPaNrrUGT/G2maysFVp9dnpEye28B4pQ8NspPybR
aEQWQhSn3QyI0SzYvBe/4R+ji84x5X1rvGuavmTFBUhvf5cEpnInfAF0FOmgd4Oa
3IXuICplihWb8rqXCIgeV+n38sz1862YSkED0igJdhZuO6PpxNp79UWd8prMz01j
YpBOZ58GjPyhuR96BcpXfaFhd1wmt6RlSny2f92NXR5xzBbyFP6rDZza30qwyKcU
57USjYHitESCnVCbdhcpvJV8T78Ar8n1/6D9wJl/7I8AwEMKvddJ4ckw5ZsgF46e
K0HhowfVwoq/QTl82nuhM9CnCns/N3lpCMrXBYJkG52WQQrKQ8p8xYGL1YxeQMia
Dx7ZxxfeSx6XJbjdL+LLEfuUdfNjb30JWwQPCDjo2aOBRLpySCX4PspELcCA+Lov
0KCZBZWVcIz7vE4dajr4OD1xIPKSJ8OuIoU2JI+IqR1HERRZm7kaWwuz+ghjVtlA
/R0Qyhmn0kylzkrQbmQ3XCPn3q7PqSDjnf01hSmgvNmGlOGe1CjShBlhBSRpW1Al
xndbkRnRdSgEQzCkN6RgOHUBHNmdUy18mNPeo14T6XDJr1/tBkF5l5PNw5BF8Gqj
ilFUNXA8T7nGXpw3dtSeoiXVS7VQJQ4mfvhZNiD1EHDq61pRkI5NINdXtYNpJdUg
X5moR0iSV98zlBLtDas4Wl57WtIg9qI4PXPp85MY321vmH5oMgdAIwwsk6py5qxP
dKWT69eMzimiWJKphwnzpZReO9gsPK9xtQlhuWipu0QnwrByDIbvYd53VbnzgQoS
5FwN8UdvfpopLSD+VHc0017LhL6wbvnyzKqlSoTDORba2mIuCptQ19BXxETU3rMl
KD+Za4Szu0RjZTdXNfDsQv7g+JqiJWVRQL9yUOGjIXCVkNQZ18MzHfarhXcaQScX
W2BuwLVBu7INnU9k0Ve3waNXvX2/v7idJJEjeadkGU8HRSUcD/hxEhB0Xxsk2nl9
l9vqdXlsnU/Yh4LvBDYzBFkk1IlcHCCDFO3IhzsTQN2RGZuOq/3pGbL+GQx29SaX
dOFRdF+TuTgh4L4tQYBKeC7nb0QsymOBPsub53sD+DTcmEHJudueI/sXSPnimMde
EmBKkL4l4+9dcXjrnufhQs0ohm/kyfC50w8OsBPtV/AYPRsSU9tylCr0t5WQAua9
2gnH3zSgZCXA163RMOxDA4Xwl1RqS/O08lxhEvJr2TMBYOSJ4Uon50ufxJTvQj7L
CojGFr3wtRI/qOIsrZ/zdCzb9am/vBh6nAUMxLzDinSUJHnE/jRH8MJgOjmAw/oR
Z/rE4SF+C68gXByKbik0SLUC9j73VQb3oXZeOWdBO5cR8MIT8qS2Sz7sqV9OfRig
yazxpRRVO0IEy02qalFIVvV/6ZPWo5WK+LkMVJdjww4tCWln7BZ/LTc9EUoE3yty
wlKig3C7By3v2vr441feKbvkBF5eyepHXAUEhqC58xeKZN37/UFi1DEhcnqOvY3/
rKX0xjYWjXxdouI8I26DZUlUTlHs7ebdtffugihXD3/yiDX/hyvNFjB0F0W3VhjQ
VubD8kQ6758/oPM3zpWTmPhYJtlWeMnq9MTuaXChS5uwcHzNNQeliTEmS5l3xL+d
M011psu7kgZwJZIBhO8e0/A4LwBN+3FUrlRzfzg6nK1ysDOWEA39opWEnREXA92Y
2KQWuRo+fWsk7MJYCwltAIXfMLLa4kbLtnt91tcNj6wkBmWW7vUL6Zpu07mdL8v+
w2/JJvAo9ScRcJ0/eBMofcfv8d2EDaFyfs9rGP1QCyV6JGv6rY4gpsBoOi9q/Tgi
o3C8Q3/L31mBdU7uHV+0v7WWYgG377K/p65vRfWV3VZRQ58WsRtxfYYy9Uaut8Q5
KHoQHSPEiWli9YTy4DBEdsvdRLjqh6+s0r/Daa2v9QvCT5XEoGOTdSgnpvXn6mhq
Ivz4aDen1cDQxBDYCjz/7bkTyy9hH05DUhGme6FGj6QUcT18kb1D0UmPy71oPe8Q
2Hze3YRYj/UpA9nCS/m8PnoAmmIc3LVyhal/Q9fmBf84jbteVLd8EbVzGMj37YV1
doWqJudpDS58cxh/JE5xckHq+Kp005+cg39pID4YE8CGEjWXZMwOpsbPAqzP7PQ7
efJg0hq008AeQT2mDV157m0aNqJh2+JzJOwLacwdQsUpWIvdIDwxzgXLObZEwoPr
JTMJ/QkgKYzPXdBh+PRPr9Uf2MpBnCTloqFNfiGOG0DwzmUabuzGlTR7XlTtHfRE
4kdjlYrGTlwN9za23772uQKDwjykNCLIR+QZt/nZG9QOoiQncSeFsZBYzpX/AcIu
Zww++yBvJmDtSeQxIJapXv7Tsp3dpKaokq4eSWT+jAz+D9DEosEAZjs7sFnf56so
OnmMSbeKCmZrZZ/hOt0rT74Y3nq/Nl9M/PyVYIJj2kvNgTo5ogRuhZ1ruEWRiKmh
Pzt9RH534M3X1Tf1BNoApQM/J8pNiu9zbInFslFZDrI6Y3SOpaotGzQ1k+lonr2N
p449zx4bQiBkG1D+DOqOR7uH2dUFKEEM0a4CbP4vDrS1j6LtgaRFQTaW38zlz0io
9prsrKyQDoILGXVRzZGlAcLnCLHXkjtbKpLqDhdlkiBF0bWQTtKs807br8UJ69e/
9CGWA1aOwuzA1yUu6GN1qi2GwrhyyDrMNDXuMh1IdxC4t6CQdH++WL9eIV0hPGx8
0OWlLP5+9WFDgWaW552PFC3zKigeclxqEj7OyanMnMlAoampc6fnczwQ/Hmh746U
dkGrfMHFES/rdZn9D5fm4iaP2giSrbyLzlTfDPPnlB2vkgvvlr93pKGR/9korPZ0
IS884ifj04QBvGWKqbosDUmYsL7oj9Jb2le6/Is1cd82JpwygNHAgvBsjjF4YT3Q
4RvNXisHZ/F61qLzMiDqmUYNTjzB2s2/PcLEsNlFdU4sFMCvCSBGsD4mcqAz7EOB
Heihkipz0t35ncn6Q6H5jKwOroCMxt3Bq+ikhu2iL1waYuWCtQIMQQpPrFZEsVk9
s4Kyldj96aInXPJ8LyXsoeOF9gOITNq60bI120W00mdIRG/sLoNliJA3UlK8/0uI
vY7HzL6djt3qdtINzYel4QMxsbhe72F06+PVdLC1EmdzixvTTW1uuCCNIlNs1p1h
utIGeJl8pv7iTH5TkPrY9rEHxYMCY6ClF3TVbu9plzhJ0ubAOlkBqS6toRITHRVS
IoKS3O2wmxKYxpU2lFNYqPeNeHf0s0bsvOQIpCqsx7IEYIIROWaiMJdSE8f5JXcw
J5bmODlMsvfIfiloSwXqUUdSBNhluLvgvTPGPKFmdJWVTdwrZcXI7tE8oms/wigC
HhcaHApkv91jo2vY1viu6NfIDt9Igr5XB1Ox3gKe7JSnEFX9Ql2bnK3IJM10KC+K
dCZ0cTh2L4KMTQzH992A+b988NZkj6+vsRRIoO5p5qddsdohLbc86AhI5sxhUFks
0H1H2fF506qRTNXByj87itD7eECIW1DRNixWU/estKuUpnwIn0GW10QXGiwxxwig
uZrvy9LegvdjmYl/ZGG9rxCsqJ1sUCls1gQkoIs3+7Ull/m8n+zbCjyxgg42x3N0
Cj5wW7mMmhZROAbpOc57F6PS8SyyA6TeCAlL5talBdC5pgGeHnKL4kNzRSW2qh18
K3b/9ICy9PZYxvOnwP0XcBFL8KN8TUfUrMJwh2eH1aJuQ81cq8/hqWOI/Kass6u+
QF/q6jjQ7KsIBFACnhExJWD8wa/cNUIidLFcIcpPQnqD9BrrncZ0p+LEBWKYkC+d
2TMG1QYMhkBZgBBpIZPq+MenaXMx5XYaiDjQwqb11hBwSc09fKncA0mHFXiRPQrC
aXlIOqacLNDA03opakUVbt3vPsH5YUo1zVeI83QYKWN0K2By5SxvlFn+oQfolkJl
7mAeY3WShUE3qgKVsm2DRCwRsAfdnw9eIC4DZ2SvRMkpRcXB+ioALP9RatBvnmhl
EraN+Q8hRRtiJ0ofGbAGzPBvXuTL+DoEH9mUkzvAk39ep1Z/qAXMB/iuTz0qVNoM
Cl8qlCru/jNzyjsVfyXm08T6dumE98zzm3wxla91EQ8sB7VT1alEDVvAFvODblIF
Gwi71Z9YHSjlBo7IRs+DwRaU+QU6LZoiBiqIBdr5SC/gJs3JD8+wfW2JBulgGVI3
kmhI67n7DvaYLlnCwcc4mVGzRpG3sNcjvqzX/jAImnW7sGvq7t37zxkAy80f98Ab
9jlpPJAniL9FLDJ4he6Ifikr42dN0Rbp839DVYBeg/43Ln15gd3XMuXkiaoKtSwq
Ot2JxgtKM9JiA6yWwu4UjvuUkarIEZOxqOHDkRO6YKNtMZ7EfCGepH/5tcPyiy6z
Lk4XoGT0Sux7EnofAmhb+hhxxa1vtKv35IpznIAB2+/JsXb92bWa+X8//CPK8dZg
qWO2SAghtcJ1ftSYjN+Zk89JMntNlPf0elqd7F9Q16d3im5GsFPwqCLQ1QXTrW2A
AuUk9aL1abROKRA46wvNkasac160K+46gpLA8EOBeFkOUrt7B5Hp5ZpOxqLgc1Hb
pwaLJxqoaGskgbVn2l/V1oip7otkLPqaeDGJ8nLAoyQbBmt0zTFR4Ir/UPIMorVX
8DhYxbJ/73jchfyng0QsJQdQNcIwv3NDPSYzQa33hKxGAsgAr88H5D+km/6/N3oe
7w+8e/GYW/DAy1b9lxGwaaWVeUT4Qyb7LArmc9zDxNRLFUQdKGb/HLnQan1DdSV0
WAjrFZMie8/IiksRcpFkk/21OPfaADqq8IquYGsdYzwAchXfSTnlLZ5d6nQcLwtK
DptrQcLzz7eTtS9usmkbq+eJH7RZ7ulKZgGDxKXMmXRJWYkUUf9i4w4dYqdVWImy
Tmd4lcvihOqQOF7yPTuqe9aNaBdN5UeJNeaQWteJaLupu3hdef8w5dsFZZovdDSs
NJB/eRCb9EYovt433VT+wKBBeAhCOASKLt7VQKLeko9wZU8uUiJ6KQAFT/ZOCEsH
mvL15IF5Ch6E6tGna1KHHTWRg34cZTs7hXiJ1oGBDC7vAkjfm8i5WJx1HaLWZlL8
PbH0id7cmJtQUhjzemBZfNYCX25BNwu/5Yh0P4ghaIRfnkY7DcmnAd+TO+dIvkln
SbwHUjJxdWISTX3rfAmtDXi6lLNJa8/e2GXHjMUDD0BVknYrZ5JEGiiRj4OrawYH
DG2khrvs9sv/AVcVoNz3d+6R0gRQrnhxFQMguaXdGfVaiX0esQDtiC0E0DjJxeG/
3s026UYfm8YuRo9GjU8aLjAXOTZ+e4b7RTyirAUoMq0pNkWyRvdmZc3wg5S+z85+
e2CEf85MyLRS8SE2Chham3Z5/M1Fc8/WCEuL0ry9rOQ/z/XnY1K1sTSox9VbKgA/
6iXf2MPswzZ2tpe1Czy6lAA1Av4/O7UczOx3GPSh64heHTvbAe0zM7Pi6Zm+m2BU
3ohm2BZtYc1HYCdrEVEtuM9MQ8HBgGueTcGFuDWwpx4da1Dn3aJ9RWhfB0RqOYKj
TypTpK35Lx0vttLWhYRZSHp5D5GRxEXnBt29VPZY4wMNk7LzQHDFxFKXTmHy6nLW
lLDODgYgYfef2SPttau/wDSeh7xjcCGp7riW9qtjKtYipueLwuwI2ZRtR9IheCaf
z2+4uzu5b6zTzgtty9FN3SijVI1W2fNuDWoA9+L/TmgjJlKz0JY0EYu5x589sb2I
Xoh4r3Lga0nvmgehvQVWByaY512dXV/EZOxMwS8QmCYozjWn0A262S8b8r2szDCG
CBXsKqvHtqx6dmp9MNjthu9o2CLMaaDzeYEZ1dT0DZhL8bH+W7D3czgLJoguDXSw
PSTYpuIymShAvgVZl/2NCzLsszmVEN4J4TetQMvS5xIz4pT8lvzeMQgcXvIFLBge
aSVJ7/D0kFfnD8o/o1cCGgbINupx6OmECLkOAPQEyvqlX1W2znIdE1e7V7fWcWaT
0EDX1I/3m6RIwHTD462PmIukPUVDJALsGwE0vWkwmk0NwjvJrdApXPxr8VjawFjR
PvJEX1ZCdp/0F2cFk5MxuWCirlNb5CZ+gB0j0tfpBS27wQoVUrkbOHLsbJ/r7Tjm
4IxWm5I7GIoig0hUpsqpvpicBoZx5ebGnMOGAw1UQDKzNYCiNCJ8SwRf1ZWxAX4M
TJiNbltfgKdGj2gRCXSm6Ja+B5Q5NDnkxmQdL/ZzlPL+4920fNZ6EYvI7lO+7j+m
vfnf65qcqXGD8wtz1NnHtSfD0aTO6ceYLHkRn6cOZ8yk20hHZWcfBbIlk6XoCWWa
TRMEQBXgI8drb2f2nRIVH7YW5Efkw/uuQa9pxSmQQHsfuAOwQvY6m/3Ho+ZMUTuY
uc/mEb6KVT+x4KnK1KthvqZvwz2J8OrUREpX5Z7XESuJstZ9uYIygiq4Dt7kKITu
KkqsDiA6sjp7BMhPGrs3hPc9bPgtv9+fHdBZKCgpc/sg1kguSk1NQJLsJvyKAJ5D
Hxf85HW+U19yjkF4dhJJkDjZGBoEM3tBV+p7gjqIUP3D4PHPCHFXQ5J73TIHklvu
qUsR0BIpt4yvF+mhvgWxqmlRIESDOK5Jt3Un+IUadfYpnvO1xN3qzr6k2BzcSSjL
ID/0jyyjTJTJgY9WCtkQcegFR3lcsRmI6kTyh+g9kwqDU7mgJa/zXYSLXS2gWRvU
1yYP2Q8YR62meh2dMgF6eEjo0AL4nGBd6ps9ZgOALEYAdLkVs96cSeuoEtqa3jwW
Fu5wAViBRqT1Ki08fF5t2hm/yDOfDVI85eJnYvq2ngOneXQiCuuoK9Wrk3++3dI1
abIxUykgfWQDhAxYpWMrP19CLj/BrjZn50O11UdxJH8sZf58OKC53hy7yc58N2xl
KScgvN6f9nN4Vjvo3PFb738LTp2LAGt9wTdKaOmQMbuOT9kvtM3AKDKnHKAcU9P2
MkpwDvBw+btC/nqnUci3sJ3XEfCongVxS8wvNLU7XvZ0g4giJtuMnq0lfcw+nMkn
wsrcPm5wn+Ivd6jxQooEND2vEjNxI3IyJZIEWbWCnUwwTLboxTPvZSOLE6JU7UNR
Nvhh1Sjk+TvQ/krgMCdFc097U+ohDY072E6JccFChUnYlyJEOT+nMFyHBdR1SXuh
phQj7jwBi3Ic8kfRKkjPKIhOsopkTZi7qT9aQil4JN30tok94bz78HahmAc7PG/w
g5CjZ4rVyORg0y1NKRrNBhAE7pVzyl+JfU36iuYt3OtdrlcE3oJoZmPfaze2DZJa
XXqrMvspbw3e31r1gQ2mzUV0ykmOfWDJZCMhZLjeBvGqjBNT0nBx620Oaz/HODxQ
cHWJ9UUen/VsnaS8k+kxWbS7ROeveaMh0iqt7gU//u/GhOYifQjL48ZHTckssY/l
pXZN90utYJZiPqbk3hqvSeUYk2cO8poauGFTYJckZvvFIerpRDS97liAGYepMc+G
mpoY2kBVulHU0rtYVllXsHlzKll3/zG2uuH4OfK8ng4NuFWAqrvT20HGMuYsCPJS
z0sFwhlLC1Xsd/u3HUT932CRUfrRRIT/Vj5melgjOX5VmKf5Z2NCzDATFVJt99Oj
XaxsRwNnKnKOB03sUJ/fYiixc2QIipssR1F1YrW2j831/OqhCYPX4l4nC8iCwzif
nCg3X9k0kWj6riRfzIglPbQaMSyOwVcOAcwnSStmfyCSefhKD6OsZ2wv9O6YRU0e
MnaxAj1Wbiheviv/7DuLamHVJK5gA1wejeXwi3qyPjbwmrMei75nbomoIS1kcQml
Huh/RxI/j289RIkzLneIfYTE0l3M/1ThnnxBqYBJEBbij8vFQ4ZUdX0DAioWjr0q
v2hwQNtHrsLE6x0FruwstQtG2KQs1HO8sIU7nqkc5ceptpM3gixayfxVTEoCaovp
5qY0yeHLK6MED8h2ZQDWdDHfvPG/Wie+7mkFzLDRneXVBvP0fj6f3seELJCheCC6
2gsCt8RqWS//JVkVurfuuUNnmjv4kQ2XmMR8FZp/4Lf/kkaU3bLGRM91+JuxyDAJ
eS4C/pCbBDkNvOGkpIV+gng8wDZgjr3TTE9a1tD/cGFAqeqWd4cN1AILyAdLNy3x
1xm6sVBKT2SSQx4wlsJv2QiUHfk951f2QnB1Jfh3TqMJ2SQY4gkOEhLJ4WZ4ZcEU
O7LIrjrxzUbJ26a37hKxihB9tZIfmMPFXfyTtxbok8xs7lEzHhPauQL+WcVjatvG
ollMhsXZgwQU8E0A3NxuorJnOGXrWg6tHPVF/3SjD6SSziEdDYYsGXkrlq3+p6A/
r93Q9A2N1eSd179v6J4/idZ3pMdM3IAmB8HZ9tTDK9694wPepQTKkgfgKE2kn7Nn
jmvk1xPpvnRhjYkYWAY6aNS0OBCiqRSLzx9lRDwyDVyTRtAJA7N0ObNFBfmIQitG
I+AEvwyi3sX61E3cp3HU17wMYBVBoD9/ZCIoeMYd9+qvhBRl7MneG5UpxawSFLhR
ldqcN32qYuk1L4Jy7TBZozHiWN5nons5d99JJ9U6OyAV21LbV1g8LKtb6Fve9ID6
bkNq3DtnKr8VGP18YH6oW0cWVC1Ufk0UOukWO27YYsIU41sgn553mTCHJEJQ3JcB
UJiDVURfjmViWCSy4UQedyGmc6OhbbZ0WF5lnHC22idKIBD2uv021dAzN0Kryzuc
ymL5Gk5oyM5cZUqR/Fdf6nYeFubPCrbEs7Fp7eGB3eJA3wPpM2//Xkwf8UeoR0ro
HHNVvzAzTPzhIHLLNYUyw7pWVSNGFyK3yu+ct3wsYnUuznp5alA6vRW5x++wSLN7
jOI3pRBCC0uchXyomnXKDV6xyfpUbN41uFLiaDt5icgzhrPJzcyjDOaTlkBR/Xei
No/NXeCAsBVLlaIpShAYysNyDvtuU/Kinl/F41OxqJnAXit4d+9y05Ow2GYFxgII
d7ZGKlmU+WMe8c4aFThD5i+w9lc3zq0+eu4ZxLE42ucgrmi6YKjJvHshj3MtSp4q
6ZBRnOBtaP9i/ScR6dJ2W0+txGIC36EHpoFbxZeR3JE5IhyrQsyxBHuvDfu0xj9I
msHEDNr9g7nIu6hZRslYnhDXwt98QwtGj1U9RHkEjVWao8BaR7+mNI6POwGYQ8KZ
JdolEH4Tux+ZI8iiUcj6tL4bGMDwL7QuuB9hQ8UEuhqKhFaxjOfRdKcNit6/Lq+I
2DXzf7iL2ctO+5wJTOQFO9/EeW5w1AInOR7bZcc/wg6HcfkBp1HdrBi/4RJ7qZHC
QYWtz/088XDQJNsxW7KMuy+pXDkmIgLFDRXYjZVJzXL/a31kbp8UnG9MBXgnyIZO
VYSW3zL8bQB9oXLopRyqFzN4aUIneu1OEONOyHWV7o+t43QD8xh6j3IieAzqCTeg
uhJRpIZJi4peMhzDFF96uiFZslK8bKurmAIUqbKj/8w4gxdUFKrxtaT0hag/gOt3
9vxud3WIopJHJrMLIpXlhvTM0V+WN93+tx5uDG0Q1B0fdi9F6Z8hJGn5pkaZg2hl
jlhplhatjjkD5Q2vgeMYVYu3uj+saf9XSPNUujzWioFTnMSyZrvfz1iESMOjPVSa
wU2KSMJ4DLffjm78uHUabrweggr3++CytWWfVP/4GfDOWra0GKody3xtdM2j3IxR
wL5v5/HlTimQQc3OZKO6ER6PL9zYnLy+XEN4cjosz4N5vfkulaY7pcAcN3RN5U9s
0avcwlxEKvLAa0gm3vqEyhP3kzQDzDNMeVNy980Fo0dI3VpU1FdsglsT6+m3tV9F
8SbqRurBr1mbRQdc7Vrb99MaSaPz5IRFm/ADOLROb/E2hVhAqq8i5CariRt09upE
VSsWirjj1pTkzDEAd2sPDW+4ETG4h6qduBSi7uoC2ytGwNb5fZkAjdhNwzsZtXvC
D3zu1BhEZ0v4IsIE8qph5nWj+2ut9Q/JV3kwvjvTj0CNGOpb/r1gJSQf2nfwfvpJ
nguXQmSkPEuDNnINZpk2bHFynXgKG6INVco7t0cQ3HDp5k55qWMsJLyoxpBzzo1B
ibTNbfW+Nt5nW5mlAWisULQHOuveQQ3DlxO6P24cRYQc6xYsOE3LU3U2fAmlKQhO
8z6iJks9DPIfQrtpDyZLhoFZGWRAlkeGnqDP7oPVsH2chmoZnkejc7SsnqdVTrQa
buTXlxdDIHqbeu0MsYFH9UtyL77mZ9O8UIrEpqAK19Gn52/0c7jeto27QbOLcH+F
QrhOYqxnLsw5z7+w02ywxrOEXHLs9BkcNWDztMMujdf1msWgameRU6jcqO0EqlmT
ZJilrbDksz5xdwZehTrT+uSNFurqha7lcYl4SHifsHPvDgY16wbf2osD7PuczgIG
xFMljMW8EJcQ2d1XdsmoUrYd68Rz41RHjBTckbNQvIJrHH35Lzznb3PrSnFzD/+w
RxXrga4KsxH+jggcYz3QG6hHOxveSCYTK5ZsPLdqhQGAQN7txhpzyckMJYQlC5Cx
Midc4XR4TSNeY16olNkKM9L+bgK/QBDU8gL802qqRktHHiPu2oInBYq8mzFJSxP6
uVFlBlQAdJwmhrKwnKz/YX5pONCeO8b51Y/iyE3M+MsWgbWYHiby7DnL3s5OHFX6
wFnHqjooQaM+RuDiklFLThIvKK0l/NetkOqGyIqJLXIeb4dJRSUISrCosLWTUQfh
qATKGPOjtTQ/6HfxaDBAWf4zYUkEidnKugwGU6ojlAaM5JhlPd6uJLigLKM/sQz3
vl9WHvUHcu6LBbP9FrfXvWuOdk5dtoKSB9rbYaTr6F6dt85g1aQshGcn7A1T36ZA
DR4utXAtajIIZC0okVlJA/lqo6XjoCOAvZSAPb9JJUVonzv3lHYiYC5WShos0E9L
guBqgQ4aRHzLZaIrNED2y/xIF4gX2waDlVIOAzcptAci6U47Dlx3qLEFP1mFOcS5
MRTJXegb//tDsDmop7MrYV8jXxCLwHxt+q8qrvD+d6xSqSkIoLzguwITrOHnkjhD
c8i3iSrOSdEWG0dA8bsP89TJHi2Du8/bqRCrsLj01LleSN0QR6Ezyu09dVkKgw4o
GQ8+rZvNwnhx3nebo5tQ2e00FNR5igqe4ZB/EEJItUDbt/CKlyFn/mspKohK546c
9ppZwF591eevjTlBgnqVI7Bsd4qCja2BPJ2Q4PTdp3YJoFWOWrRWmN04NR0c1RSN
qPMCDm4qaclCXtnwf1XhP94qnHAm7wmjZGJNG63cAnH5tpwLuQ8cauS3Sz7zy7/F
RhytLKemOsvpsGmGmWTSvlwSbj2k5D2QRu6i6mFIFdVrEGE5C4Dsu9/is3LyaiTd
b6zeVP7f8Pd55oTu5r7no4tapbdayEtuLf4l4txV08lspZahG1EtbDifk4bH5jsU
hRR8SdmtOCAe9mIhFTA2F9qTcSIB9rA8FNSn1DNfQfqE4Q3+cceyf0mRD8hVYux7
5MRfB81XIPfAR73izcbj5OHN7xAjvso1tirErW5lEmG99hchDw6lHLKZ/p9zubMT
6kjcf995EEmNsYxkK5+Knq+13rHRIna/a+SIWH3U+PH0PwEbgRz+wZxMOU9uPJUO
+5wZLSlvuATiyt8wrpJ0jObsaOVjjSIh6hqgbkCKR+PHqpGkLzI5jGgsgov6kAmA
tnkNVQa8WoDNyws0JjmTuGBJtnUJ/e+583o1qPA6bKhpLBfg4uhVRSEZ1YkL4U+7
l9zeb9q30o6/+F2Z0WSOw3srIi2ZBUpsdmXKLsIS1dVX1bmxLx8MthWTth5hIj94
eatCeLnNu/MwAQ8xm4t3cEzT0SvpDsYB1fzUjPZyxa5rHTaed5G1c089v118OK6m
t9CkWXP+IzF93Uplwu+QYsfbULF3wMs2VW+ZjgfqfpdzOVjIfaff6vyM+ADJeHYl
7q3djUn2JaKTC3nOFbCCIgWs46ZAiPI3+0XiixQp4YbY05m5nWYdnU8wITEE2KUS
hpPdXedItt8Iin7iP97TY8NpnPTQCun3BqyFC7a4qGrN/H+ZkCQD85QL5vdpcLY/
36xRsX/BYNePigX75W//Xqek41gqwKbcp3KnxKIh7NujEZhCPR0PrgCLdYg3s2xX
p8X7wnVW1IV6Ihj2ZCi9r4x2upDgUrXZZwLp/FfbatSSA1SGxPgrm/KEErJ21AOR
Nn5lAlsUNiHvXkWt6D7Hct97hXc3DyKUf7zgXIKDXcjpkMR4G1AOEh5ZVdTMiCxu
33B904cd7dqHA12GdgUxrsQVETsjFL4dNS/FmO5vyioZXvCYC3wXQyV8j2yAuvT7
us4ZFV/d6ZMGztROjtHIytJ2r3mPBkSFdQk78qn51fqI4Lns1kMRS2GkC48pK0jy
7gehw54OOpfXfF0Wnc/F89qNgx+NadEe4NtOx/Sc6EOEj9b8DVxd/9mMQWAnYyjt
irb47iOkOtVYw27ZmUKtRMdwkTZTxNJK65JT25S8bPMh6t6ooqovqH68UihdBhT0
cymbilaeTcfbvmaUXudelPQvHHfTfqPzd0wzPgtjh0mzMsIUZ8jK0IC/ALs/1+yP
/IFOmK6+tyF+JObPleeVH05UgUK7/uLk/tVoRK9L7cZeakujeOlFqAWR7wMiLWjb
gA4r8D7Zsh5AnT+SzReR+FRBLpfk/u8AF5SQeB1ohAGG+cAJxzYXH+qYZGaIsiJA
PRFc5ARSa+l0avNJ3U2ecjDl9TnKdWMYJVRW1cP7YENpe1stO/Fj7o0ckuZRE9Qk
dWLxxVrQcltZRqT2QXIfOnw/mIkK/z4DUEFTMEzVl4eoUwCaZwcE10WJvqO/QagP
okgpgnrWnVwvq4bYVMH+Y/Uq0cJyvV5g/ctnD12jg0yBFXnKEWXBPg45BLGJTNsB
7mYGPrt5BQb8EOYSmE2RnKu32nn2B3Bsi8moZTHyDiaG+6xtxFg8nvQ+Om+sJLPt
BGuDgQMzoC35INHMrNK3IexIk+3ekC8kSmmk10jSbPJZwYmuUk8oJc6B9OA+fSuw
2pF7Wg/WZoTtDrxJFgA5iuMVCH4l1dOpWB7GmldgChZpMH24Vpv8LTorO6l8Tfyu
cqgFOudbt295EX4xhTVfuanoJcTlgJAIar+CGEsk1CI+TiDr6EJFKQ+z5XOiucl9
2idTPQI0r1n91K71hwtPQjVy7s/MMSH0Xd/QLph/6HeVrQPHkJA1MixsRqpnq9xT
ck59po+DOrH8E+jReZjyE3V/1kTCDjVZsndxdizb7ZYvjchQRvtJDPuHtblKhTY+
NEZmRex5XUWvbnkkJ05e6D4evbxzSLbhB+avOzkcXIeJDQlbqvx+tjuKkuuby7TB
1C4gTyUauF0h/ddZsA7NOXRc0z96lRgFWCBRxjvqpaJfXhl3/tAene2ix+BsWH7t
+byXIlfVgauAKrnBfPzdMgosLnuPfK7v1hwwfRiZnEetgaGNUBG5VJGF8esLHyHl
k+baf3u7qh4YJb2pm3ycH9VY83OBuiKLc7BRzHV1iqAmxTz7cPhpd/Fb/sd5pTWy
8/m/blHjAnNSI9IOPxd+XfJyWF3oaPjeEBvwI29ZmW/5PUxelLzXYYAtAB/kG003
tFipFgkEZPZgnfMRZ+QJsUZeExUNT63OOthRsqMJKzLNz8QRv4hSruJD80xKpRlq
do2H6nskqfxqNvAfmQnzrkB8D4VuqsXeGa6rMuBgr2JfPjxOoy7ytBK67YYiFBOu
+HZxbZVfp7ybZIWTwj5TXWsOXj/nTdJb7XL75TevkVVXolalx6eEZW5/gS3NJHea
bA3A82oysJ/f9ayDIVM1VGGJoCZiKJJ17On1OvVm8ufjpl0CfZnOaCNqLvrn9aK3
caRnhIoG0jhIAYBZBWNCWUjnuJw4+v1UUtrXK+hWut9hjtSw3F0GCXru+TZYU3a7
zFqwjFvwSVHU9iGHhZHPUfYckgwuYcEqk8JpSAA4sua0xqsmR8IOvgZantxZ2shq
Z3EgwAuBpuhWUBG9QMPMWYfZQMONhCUudGEJ6+CqovtNrqI574Uek4nUiHRxrzjg
aE47+p1lZoq1d4E96kRL6TrLC2jaPnPDuztzDy1DXjml1QzOYHs4D5Y5PIKfrHOT
O/vmzi1QmS9SQBG/DSqJGa8hVXADUoOG5hCGByvLujzq62SMDG0zIQjC/0FGu1xh
NNStqvvmz3sCJSCH6w/mQeRwrLB5/KttClIMqTW0VzyfIYWtch8cRwxuyn2B9d3x
tUmvGzFAv1gOZ9yigVyGyJU+xhamCvwiKgI8rQI03dQs/CUokdd5qNbtrgCnfW07
MdXj0+HVZbYw0wm1/EPEVaFZH2wCDuEtYCKnwS1/wnld6t3aPqrEn460puKHqZoo
vELV9lDLRuewcDt/JVZGa+8ysSjpv/OmN5wzL8qz7H7I7xPZ6S6/XnzD+vvBtSio
aTLD3H2cUxBzY48AXdmfd/YQB8K2kRtt97a1r49qrUW3nrHY8SD005FhPg6TsJ7T
Tw8bgjVeHRSJpXdQo+GS3uhXiEpDyGCYNnNxsLtDVyuQaVHo/iuaYZqRHKK+y0RJ
uAFQ+iplxcXKLjVLm8oHEB2G+VkWNMQ0qQwTjf8U5xgUfD3jpmn2jKnamcWDUVXJ
vJsncurbp0qeRdgkdVMTCIFZoFR+jmm+dmAsYJpuebEGOwpskDDqZlTD7aZxSChs
FAR8rAhRAQXhRUmoQe7OvHAaAKu4zV17oKfmAEEnnvHq/4B5LjLiL9UQVGLKl9va
AobYktJSgFAWyM+TGtBgt0GXylugE7IggGrF6qhRSU+EJdAoIiMXaybcRZT1ztvl
IzndOaf6gM1muB9NvoRhYFrwPrzs4oPvLtDnPCD3Q02FR2FzSv6fhaL1G0G2GMmN
mnI1cYvbA/lhyALczi7HQpxt17nOM5C2h3lEQJQcbb2e53HMzFF4dtUG+2J6Nnc4
FXgFJ9jryQHbpjmhjiOGXEwMn7rCvpZIDMg1EIoSRVYs4QAPOFtrC1rBmcUHmKTr
9iQtA6uG9Dpz2v29YDbRXU30bjLLA6L9bQh66ibaxbk8xvJAVICHH3Hl3wnz+hOj
OTgCZ76YDBQ6rbi3K8iHuITeWipDNGVvf+i20mb36FPsAcl3jydjNMblVY97kkyL
y9iCo+5tOuf4BfdpLnmoTqm3TOvirVppjA1dBxQOtuyVbrBEWFZkcIIfjOcn/flC
Br+D6PZrt2Vz0CTyaFcJ0pDNXN2BCU80y7qCDDJ3Igm3NBdDJGrBsJS7SkX5QKyd
2LfDnui1tu2gdcALWLv0sliwbK6eAOq9XRlaDT59uN0dGx7EdnBluoYJC/imkIkp
AnpDHPsX9daTq6u8Owmqbtzc7p6frI5WjqN+TXV09NP5T0uPrzPoO0ipIGow/eZT
G5xC/s931Co1hFsxd+jQP0ToqVu+SRy+6rkHx6UsGqRmyHLiIKE/khe4P+9WNM0/
xU0xNz77qbY3FgcwFFOjRuCYLBiGKD0zbLXEwUcj61Tuw//9qN3k9bO7JBzyrKV8
3dfvBT3sMY7tUTX0YVXGPGd2NviCB8ClOk0EZgMbH0+jgFA68ppUZv1LWvo/aF24
0uGXsYeCClJlD1BYZkZYWRQdAQnPEaIIXnwVhd4LKep61t5Wq/BnheQwFyryl+hp
1Ptl67nLQSoiOGMBEDwhpOzOUuu04n4Np9OP8uyP5n9N80QIbBW/dMysCtTvqyuj
DMBKsFOx+JXRoFtRbA4/wDeMT7Sw48KGKMuQejCryoNkXW35lcDmp/MfcuGd3xR5
wsDdC0UKeaMdtRlfIFiip/YJlOIEYBODv6guDMQsGg2QXEMJAlRDj4H0AzTIUaLK
gQc0/+uJ/J9HkMP5NXrCcelOnynPaSMALvhBsRWlHJPDmRKRRsIDVoIfd9aeAWDH
ksIEJwFKO9PNsC7noUcw9AdszOoxwSmon9aJGcwM74FYSrcY9/pjG4AqZ6JddmWH
fABRUtuqdqOCxcy54EdOCLyQwUFqMi+7BJ0gtvH8LlfLPxlaCdiv0wmuWiaC9SUR
Wu738vYv6pi6n62fLEdyRT22r+SDFDKwha9TDO6ortUk3lvYuEWmDjMPrQApFRfv
Y27LNC4DfjK5WtNmJpdzZl+EokGgdw6LSjlA+j6RnU0bjUHP0VB20hmJY7wEF6nA
0krT/y1hhC62Om1HI5BimixRZ4lfdnh7jmmC4xnqR5SUHp6oC5CQSQj1Upccw2QL
iS8SiZ+zx7CYJuPGej1qpTjCZEJXYeWvLFhHcZ3Aq7D/j3PeJYqENRFYGuremQA8
ZvB7NcNygG1hbcSU4vN07aNMGPNjmpm9lBVtglGhCpK0xxzG53Y1auDEAbgPj4BQ
m4XqLYYK2JU3IfifcX3y1cb5c9WqBAMRilKFBTXfMlYEo+gYtHQQZNkLx7qHGKeH
5rAoItAwe6SGGsdAF7yO+JpQC+6+qViFgfHQUK7YZ11NlFTE7E0hDnpNmSmxvdWg
VwWNBm+TCORkdD944Lryh4r3/KvZnsnU/dNON97xuB30PWVrzYTgBxJpbYApERO8
gL+FqP/36BlEp2jhVuUNIWx+nOCXdSqqwz/bkCb0wp1+Q3xuDbFYkPDPFDsMQpEK
7otefhtKVwu23/YaeCAe2RKhtJyi2ov+Hktpw0Ex+W3B7dmKbWB7MXs1vit8swJR
TmUBwlvrJfomBov0V7RYFdXMq6eyRr74nH8NPKRXJ1DuxAwwED8A9OZZnZ2OEByr
xVm3s3U81Mqexm85DczHY0NlQzRl2hG7j2X6b/lol2LJVCvK6rHa3QZzRLPsoCa4
haqbBvHNiYqUWumBRfTukTqiIQIwJzAANdlu1Zi+heIQxAkS+OiAbaWgFTy6XWJ5
NSG1K2i9f9DKdSu4jXEK7NXgYXugBH4BDeqifPOr1gy95yrPTMKJ71Ag9RvSDgSA
p0+yEa+1zYVgVC5QpD1kggH3Vwk1Ck5UtcaoSUxfVoABccGaSJ1XGD4maNB9ZWth
fD8RM9kcfQA16/z1feoXRMzuhZ5MIaOXRqrMFW6/ARa2ujbY/Abf5/FtU0HS/aBn
ghWKDj4Co6DUO3y3u782HJgLyJfe9x5Z2xOr72UHzlzOGwmN3Jg4riUlDdohlqym
r1RECt3YhNwGr34pcJKy6/JrpdmnDIBjsUNiX+t/d9pz+vi3tVa8mLwseiGUfI7u
Rr7D6pcJQyXS0So0i2TQSQYTqmKVmtI7Zr13bWoeHfdGI8mHzbNDVzyCKqIdiXuK
ZQHoe/ZgxW9OF9hTcyZY464iUmWMk2NuHyCS0yUdojisb25xjNJjEbfTDGwzSOI8
qnBqZ9Uc9qnP22HzAkIoGwDl/D5AuHm8uCWvb/PPiO0SDthB8L9YgDeghVO9uxS4
15AGPyCPeBtlJPAvt0/BrOyMItOTExdBcQ3ohaHa6SA5Wu57NNVJyzZFCUNaEz5N
85Zx8Ti6O8uM4JzFbZRU6Fj7FwzlwizQjG3YAeyQPb+mByBgX+leemP47wVQqzJc
VDVu1I4KXVHIK4FiaPeVuVUZ5grc3/SuhMS2fiYW5klIeYhB0hEdrrBD3hdFRTkj
0xEaEudYd6o3C2JKcefN9KkRt83OBsruzK7JaJ6UadxMK4B2xJFqEq+MtPMqBmYi
3ogLrhExMRRVfOsGqnhqmTAXOvWT537gyGdAGvIqZ/huU3jJxWi6E1Wi7nO8gcHK
zgSKVPHcXDZm7CeHM7gqEi+17OINwhMNjB6vywwgNKTrnTUfQfbeWb2p03QAfyLF
KL/XUSyuBl1j2VWJK44MEhv7v4dqBz+X9WZerRlpNl/p8cZ/SaLB5T2Y+baBIXiO
TQGgxyVBnEVPvJ3MO0jHato1b3Do+vXxUENJyWAG0H6S6fT6IhAaY8oJgnJjbn7d
vUXdvrZLJu/2ewuXkvpsI2+b9DbVn/iUbT4vpihyGoYuAMFkKq57SLr+2r8DnGxV
SlOO0phM20G4Qb2xJw1TYrSHUFTBiM2W60Agu28vNppIyDFnMRHzdcS/3NXOvxRD
x6YjOvqszFyMfUMlDnB47zQNS+X0j5EtuLFYh7M0G+U3bGKy67vrNMeK/h2FcMcR
iqg3glqpzS4VqInPX9LUt1E+FZoNWK6myOznGYs2Xgrl+hprsj1xccv3qhHNjLQb
g9JlBve3toCDmbVKP6zsCK9I3xooAtqmssJU6AJ8JUXbun5BzDJ5kFvDsuKStx+S
usgbyRyvxMEaw48wdDZa9+3jx+/QyhVU+Wk7ucRnlrMSEzVoSAE+rNj7/HInVTgH
cRs1mf4zY6e3R3SAT0HDqAuBEaJk6Yp1yYNHJvoPVUbK3S5vMlrNOn+khSFlhEzp
ILGA9CMS5f/Aaw0es0X3WsZFdElKXVMVm/Dj2UhPo6Of6rzRUjyU+yfinJ1IrWSW
Pd7T3dmaOE8ZCGtE92ud6dHRR+D8Yl9DmIB1fKtU4y/Qx5okFwoDS2LmZD6OJkZu
4t+Z5vwLLS4EByZ+TPgmRYF9a5FCuKH23qe8BOg0vhvb3Cy6Q5U1tFRb/woZIP1t
7H+BZMamHuzoDMGIOx41QQOWuUYe6a5trHZtuyR9VrVBP+tI0i1SOw7s3UcePN75
zINxZqbq/m1PXPGFxHAxrBQ1f1AE+20O5Yv+RZME90NdvLHhnm7VJjE0PdwjlT+B
RzztOvDhYztd9SoDgtjo33omwCzZ01DSvlb2qyTEk46VNPwZWxTr5OLzHlStDtSI
B7KqYsLtoMQteUcH65esQjyRp7u22Jvr1QvRMkDtrEXFGg/dGc70UFFVyzYiUrQA
/usf9IS+RF/v56HhGK1gwPfSwZnO2VyhPUyOPEIL5NLs8FzUbhWtpneYMgGQYsVv
2erbraiEgQxR1wUOFa9FW8pEusNkULmQCwCIQTrBI12jyW/66d5wjjjSjqcQyBeO
Q6iYPcze4nopbhv+D5UR3/+BteFcE50ztz+ot7HH7hHK4yeEmEcTYBw2N/wblr9v
FaEIkbbpkdL2pYgKegXDeGukmCEyA7DNDZvPQcHFBlagJirSNptLn8p+JKYG+quv
EUdK8VSThGt7AJzgQNsG6k5nurKmgWukBCzhX3evq1tyG7m0q9wyZsNE55gfb+qM
x+b4OBZbIbAhivqyPwIUoIb8xOjI/SG1n+4QfSzdoxTQdKMKMK1h+wvcHpDaOPdq
GyklT2oq3PoZomWJPdrR+PnjTDHh4HkqpCz9Jc2ZeFxzfst4agvEOqPTEwKV1urk
bB09+wNYRAn2Zqat66ZiZxuYvJLlolZIbow6PEw8tEu28JhQksBXMohBF52FsSRI
tqV6SlG5euHDpm1Cn0VfF+svTwRzs1Oi1O63kQ4vs43xn3P3jLqNwSJRQwtSSiXF
81nUf7yseDPoWNX2030CbkmJcufd/7iRzOhQ6KJJ1zf6O/Z6+QYtZQxBa1B9S1z6
ZAQtlBK6yLocRUDywWK8NjA5NfIVJU0XZ92DwGHzi2VL+ENyof82vWWqwfak5BF0
wdUB9AMFxlCcJPtygT6zEC8CIW/kwdV8DFD0CO6RSSif5Yb9lH174gXjsEBGUL1i
IEkp/nQbW70hFr01eKkKuyyqCOM8BrV/M5X+vzbpBJOSmDMgD2kiA6vQ9kQ+8f7Y
0zTi2lXTwO3GCWLiIIGS5lanIjEz4EmBYB1Liyl6l31RrQ6PAp0TGDBgcNj85+gP
4lS1KEZibOHAr6MiyEQBQDGawT7T3CHHXzPKVyv2MHF/tK1i8KS3YmhfFAbLDDnB
4DYBzGIBGc4jPLNYCJCdLFROXoHBOntKJ8iCBspeBtPUGiD4+ppdj5BD8Bm8oqZu
MhnzG2cTIJ+L2xlW/hTX/vVkvyT+M/gJbQQcZvmmRK2YMShFWEmGaiyloHa1Y7W0
rVl1bR5DunhJnKYxFtYbE7QT1BZBXwkIJxyWitde1563KubnWCbU6/1oqXuByF7w
51WuR+xeHk1Rvaj45m+hUxvjAOBngGyw1khoDm9j0qg2zROjtPtL4TPvAMTyoTFh
FLIkBRlWRLik0th9TC+kMDPWy/XrRupl3qG8kqQHrf6Z/Df6xg80oXuZyJYdaIQU
N6VE9suO68H6hoFr0Z0sNY9JMY/HqfLsSdcwMcP29lZa5wEhGyzEtdzaZwH2Iomv
Wagx3F6jX54LXaQgWp6hYRxA0C9cBTNDSMbtDmVeoTQARj3xmAcMX1AS+ff3Xozn
nDbzFI+PxcnyuxiFScZuz9EcVNH4AVSEQZuMBQy99lfVwIJq5AStW9/w2z1IFXj5
Osb80xRXPtSw0RXy05+shxQdZxRSiojK7AuigUNb0UOuYJSvda8LumcwXuurKRav
DtvWQCm468nlrPGmBxgkprYM0MsGS9HjnOE8xIAioxoGz9w+XSuNjHi32wma7iTi
tL/KP8q4rvbH4Jt8FkxxhDlfESRdOCCzqmLGSu7RuG7NawoHzNHov4iGBH6kZvRg
DQQKj7eU1gxECnTijc8U3JB4k/xOhwMdfj8Q/vU+TFraJ5kcEcatv2QmhI1xA9qI
7V8ioAthPbGruACsT1eWbDzQNpC+Q4zJY91Jx3TY7UY4Nnp6F9W+J0ASs46nm1MA
LqbBbadJZdPlm1O84z7rwd2fDK+ait5f7BQNrFUA9gVdU4g8FgbwLaKES/mq5boJ
GVAPt97dJhtNw8xT3qAFVqcl4DSOVP4XMSduqD1dR+/h6051GL9NGW0/y7X6eMmU
wQOJ0zFVY3nEWAuvauGCTMU5YID3d7K2hpQaj5BqPqwfcP+xPoQtrRy41Pq6b5Hj
u1/sqcP2YJSDzx+QFG7YH28WwaVPn7tq8T4a9CJTzinaxLcJe+5nfAtN/6i9DQ31
Z18UH+bxQrt/SUMTOpnu5+4Y5pkK4G6491+CTWNpR4AG03jbtwgB3Em4i7OvJkxh
AE9mONmiqZEaFx2dxSenbz3BgEHZIOIDSfdqgaaPuF42JlnE2mq7B2oocbaObwdX
MCBrJZgIoTlTNBcQx8gclCxU6NiMuSeO+w8ttsqj/wBMW9OBOaEZvINBicyyg3k1
JvwZ2AZpJC2mYRTUTX6q/zO/oeOVwdwQCA2Ql1pK10DaZpm7aym3O0d3rw5/uu8I
rGLmmPIWOTnVLjOR7dZUbazbzYtPprPFl88hw7viDW2yOUvpfCTLNAJWd1IQ+8TM
dNrO4K66163KjeB9bc4+TygRx/WMrVTFRxOmosO2j9h+BCw6DVB5lOAB3NoTo2Uc
P1xZT1/w8LeqXh4vAA4paihpyR72PP1T6q5D4+B4Pnfm8w6rDOQBOWPiF+KI3Azk
Zybqh3lB8OXoFttwiWaxCUddNaobVnGn8YTDt0lmN7OSrGz/iNSraB7gFRSkRdUS
RIVM4DNNTAo3NsjRUl/zdxMXxMggxYZ1BBG9jVIPJLPS7lmQALjzDGeL0yCNegwP
ml+plEQKKMHNcc/xsVmLuo6Zm6vBwLPVHMME0UYBQEnk18Nn+TGv64rUw2w3YcYX
KTjzzPiLFoT+L7J6C+B5TDKYn9dgvsKr2HWjdae2JRc3ILxzzhHB48xRFFZmo5lD
3tclxORgAZ70XbtDe6gM+3NGdGCTUib8sQfjp//+wvMtxfjj+lOnI9xzJJ6musUw
tEcGwzLMQ6m28vW0/PI7rOanIrg1VQHAkYcOSIWP3OvUfLMOZThDL2uXYmyKhSGx
GfKcKm2OwHQm78uB4XHA7rrXYPbrp/O6mKAW8K86wPVurtGHEym9YfDK6IrWD6ZK
eRcp4UE+JQ4CFFrwTafe5U63g77DH3Tzv2JOsGRjHbHw8kbHLBn7LwdHl6mzYwO6
fu+zNXRbnQF17xNNmDt5tIdaD8/QHlS0ePHmJgOglbQ=
`pragma protect end_protected
